package event_monitor_pkg is
   type n_array_t is array (natural range <>) of natural;
   type n_matrix_t is array (natural range <>) of n_array_t;
end event_monitor_pkg;

package body event_monitor_pkg is
   -- subprogram bodies here
end event_monitor_pkg;