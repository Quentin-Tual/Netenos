library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
library gtech_lib;
 
entity source_altered is
	port(
		i0 : in  std_logic;
		i1 : in  std_logic;
		i2 : in  std_logic;
		i3 : in  std_logic;
		i4 : in  std_logic;
		i5 : in  std_logic;
		i6 : in  std_logic;
		i7 : in  std_logic;
		i8 : in  std_logic;
		i9 : in  std_logic;
		i10 : in  std_logic;
		i11 : in  std_logic;
		i12 : in  std_logic;
		i13 : in  std_logic;
		i14 : in  std_logic;
		i15 : in  std_logic;
		i16 : in  std_logic;
		i17 : in  std_logic;
		i18 : in  std_logic;
		i19 : in  std_logic;
		i20 : in  std_logic;
		i21 : in  std_logic;
		i22 : in  std_logic;
		i23 : in  std_logic;
		i24 : in  std_logic;
		i25 : in  std_logic;
		i26 : in  std_logic;
		i27 : in  std_logic;
		i28 : in  std_logic;
		i29 : in  std_logic;
		i30 : in  std_logic;
		i31 : in  std_logic;
		i32 : in  std_logic;
		i33 : in  std_logic;
		i34 : in  std_logic;
		i35 : in  std_logic;
		i36 : in  std_logic;
		i37 : in  std_logic;
		i38 : in  std_logic;
		i39 : in  std_logic;
		i40 : in  std_logic;
		o0 : out std_logic;
		o1 : out std_logic;
		o2 : out std_logic;
		o3 : out std_logic;
		o4 : out std_logic;
		o5 : out std_logic;
		o6 : out std_logic;
		o7 : out std_logic;
		o8 : out std_logic;
		o9 : out std_logic;
		o10 : out std_logic;
		o11 : out std_logic;
		o12 : out std_logic;
		o13 : out std_logic;
		o14 : out std_logic;
		o15 : out std_logic;
		o16 : out std_logic;
		o17 : out std_logic;
		o18 : out std_logic;
		o19 : out std_logic;
		o20 : out std_logic;
		o21 : out std_logic;
		o22 : out std_logic;
		o23 : out std_logic;
		o24 : out std_logic;
		o25 : out std_logic;
		o26 : out std_logic;
		o27 : out std_logic;
		o28 : out std_logic;
		o29 : out std_logic;
		o30 : out std_logic;
		o31 : out std_logic;
		o32 : out std_logic;
		o33 : out std_logic;
		o34 : out std_logic;
		o35 : out std_logic;
		o36 : out std_logic;
		o37 : out std_logic;
		o38 : out std_logic;
		o39 : out std_logic;
		o40 : out std_logic;
		o41 : out std_logic;
		o42 : out std_logic;
		o43 : out std_logic;
		o44 : out std_logic;
		o45 : out std_logic;
		o46 : out std_logic;
		o47 : out std_logic;
		o48 : out std_logic;
		o49 : out std_logic;
		o50 : out std_logic;
		o51 : out std_logic;
		o52 : out std_logic;
		o53 : out std_logic;
		o54 : out std_logic;
		o55 : out std_logic;
		o56 : out std_logic;
		o57 : out std_logic;
		o58 : out std_logic;
		o59 : out std_logic;
		o60 : out std_logic;
		o61 : out std_logic;
		o62 : out std_logic;
		o63 : out std_logic;
		o64 : out std_logic;
		o65 : out std_logic;
		o66 : out std_logic;
		o67 : out std_logic;
		o68 : out std_logic;
		o69 : out std_logic;
		o70 : out std_logic;
		o71 : out std_logic;
		o72 : out std_logic
	);
end source_altered;
 
architecture netenos of source_altered is
	signal Not60_o0 : std_logic;
	signal Not80_o0 : std_logic;
	signal Not100_o0 : std_logic;
	signal Not120_o0 : std_logic;
	signal Not140_o0 : std_logic;
	signal Not160_o0 : std_logic;
	signal Not180_o0 : std_logic;
	signal Xor2200_o0 : std_logic;
	signal Nor2220_o0 : std_logic;
	signal And2240_o0 : std_logic;
	signal And2260_o0 : std_logic;
	signal Or2280_o0 : std_logic;
	signal And2300_o0 : std_logic;
	signal And2320_o0 : std_logic;
	signal And2340_o0 : std_logic;
	signal Or2360_o0 : std_logic;
	signal And2380_o0 : std_logic;
	signal And2400_o0 : std_logic;
	signal And2420_o0 : std_logic;
	signal Nor2440_o0 : std_logic;
	signal Or2460_o0 : std_logic;
	signal Or2480_o0 : std_logic;
	signal And2500_o0 : std_logic;
	signal Or2520_o0 : std_logic;
	signal Not540_o0 : std_logic;
	signal And2560_o0 : std_logic;
	signal And2580_o0 : std_logic;
	signal And2600_o0 : std_logic;
	signal Not620_o0 : std_logic;
	signal And2640_o0 : std_logic;
	signal And2660_o0 : std_logic;
	signal Or2680_o0 : std_logic;
	signal And2700_o0 : std_logic;
	signal And2720_o0 : std_logic;
	signal Or2740_o0 : std_logic;
	signal And2760_o0 : std_logic;
	signal And2780_o0 : std_logic;
	signal Or2800_o0 : std_logic;
	signal And2820_o0 : std_logic;
	signal And2840_o0 : std_logic;
	signal Or2860_o0 : std_logic;
	signal And2880_o0 : std_logic;
	signal And2900_o0 : std_logic;
	signal Or2920_o0 : std_logic;
	signal And2940_o0 : std_logic;
	signal Xor2960_o0 : std_logic;
	signal And2980_o0 : std_logic;
	signal And21000_o0 : std_logic;
	signal Or21020_o0 : std_logic;
	signal Not1040_o0 : std_logic;
	signal And21060_o0 : std_logic;
	signal Not1080_o0 : std_logic;
	signal And21100_o0 : std_logic;
	signal And21120_o0 : std_logic;
	signal Nor21140_o0 : std_logic;
	signal And21160_o0 : std_logic;
	signal And21180_o0 : std_logic;
	signal And21200_o0 : std_logic;
	signal Nor21220_o0 : std_logic;
	signal And21240_o0 : std_logic;
	signal Nor21260_o0 : std_logic;
	signal Not1280_o0 : std_logic;
	signal And21300_o0 : std_logic;
	signal And21320_o0 : std_logic;
	signal And21340_o0 : std_logic;
	signal And21360_o0 : std_logic;
	signal Or21380_o0 : std_logic;
	signal Or21400_o0 : std_logic;
	signal And21420_o0 : std_logic;
	signal And21440_o0 : std_logic;
	signal Or21460_o0 : std_logic;
	signal And21480_o0 : std_logic;
	signal Not1500_o0 : std_logic;
	signal And21520_o0 : std_logic;
	signal And21540_o0 : std_logic;
	signal Xor21560_o0 : std_logic;
	signal Or21580_o0 : std_logic;
	signal And21600_o0 : std_logic;
	signal Xor21620_o0 : std_logic;
	signal And21640_o0 : std_logic;
	signal And21660_o0 : std_logic;
	signal Or21680_o0 : std_logic;
	signal And21700_o0 : std_logic;
	signal Or21720_o0 : std_logic;
	signal And21740_o0 : std_logic;
	signal And21760_o0 : std_logic;
	signal Or21780_o0 : std_logic;
	signal And21800_o0 : std_logic;
	signal And21820_o0 : std_logic;
	signal Nor21840_o0 : std_logic;
	signal And21860_o0 : std_logic;
	signal And21880_o0 : std_logic;
	signal Or21900_o0 : std_logic;
	signal And21920_o0 : std_logic;
	signal And21940_o0 : std_logic;
	signal And21960_o0 : std_logic;
	signal Nor21980_o0 : std_logic;
	signal And22000_o0 : std_logic;
	signal And22020_o0 : std_logic;
	signal Or22040_o0 : std_logic;
	signal Nor22060_o0 : std_logic;
	signal Not2080_o0 : std_logic;
	signal And22100_o0 : std_logic;
	signal And22120_o0 : std_logic;
	signal And22140_o0 : std_logic;
	signal And22160_o0 : std_logic;
	signal Or22180_o0 : std_logic;
	signal And22200_o0 : std_logic;
	signal And22220_o0 : std_logic;
	signal And22240_o0 : std_logic;
	signal Or22260_o0 : std_logic;
	signal And22280_o0 : std_logic;
	signal And22300_o0 : std_logic;
	signal And22320_o0 : std_logic;
	signal Or22340_o0 : std_logic;
	signal And22360_o0 : std_logic;
	signal And22380_o0 : std_logic;
	signal And22400_o0 : std_logic;
	signal And22420_o0 : std_logic;
	signal Or22440_o0 : std_logic;
	signal And22460_o0 : std_logic;
	signal And22480_o0 : std_logic;
	signal And22500_o0 : std_logic;
	signal Or22520_o0 : std_logic;
	signal Or22540_o0 : std_logic;
	signal And22560_o0 : std_logic;
	signal And22580_o0 : std_logic;
	signal Nor22600_o0 : std_logic;
	signal And22620_o0 : std_logic;
	signal And22640_o0 : std_logic;
	signal And22660_o0 : std_logic;
	signal Or22680_o0 : std_logic;
	signal And22700_o0 : std_logic;
	signal Nand22720_o0 : std_logic;
	signal And22740_o0 : std_logic;
	signal And22760_o0 : std_logic;
	signal Or22780_o0 : std_logic;
	signal And22800_o0 : std_logic;
	signal And22820_o0 : std_logic;
	signal Or22840_o0 : std_logic;
	signal And22860_o0 : std_logic;
	signal And22880_o0 : std_logic;
	signal Nor22900_o0 : std_logic;
	signal And22920_o0 : std_logic;
	signal And22940_o0 : std_logic;
	signal And22960_o0 : std_logic;
	signal And22980_o0 : std_logic;
	signal Or23000_o0 : std_logic;
	signal And23020_o0 : std_logic;
	signal And23040_o0 : std_logic;
	signal And23060_o0 : std_logic;
	signal And23080_o0 : std_logic;
	signal And23100_o0 : std_logic;
	signal And23120_o0 : std_logic;
	signal And23140_o0 : std_logic;
	signal Or23160_o0 : std_logic;
	signal And23180_o0 : std_logic;
	signal Nor23200_o0 : std_logic;
	signal And23220_o0 : std_logic;
	signal And23240_o0 : std_logic;
	signal Or23260_o0 : std_logic;
	signal Nor23280_o0 : std_logic;
	signal Not3300_o0 : std_logic;
	signal Nor23320_o0 : std_logic;
	signal And23340_o0 : std_logic;
	signal And23360_o0 : std_logic;
	signal And23380_o0 : std_logic;
	signal And23400_o0 : std_logic;
	signal Or23420_o0 : std_logic;
	signal And23440_o0 : std_logic;
	signal And23460_o0 : std_logic;
	signal Or23480_o0 : std_logic;
	signal And23500_o0 : std_logic;
	signal And23520_o0 : std_logic;
	signal Nor23540_o0 : std_logic;
	signal And23560_o0 : std_logic;
	signal Or23580_o0 : std_logic;
	signal Nor23600_o0 : std_logic;
	signal And23620_o0 : std_logic;
	signal And23640_o0 : std_logic;
	signal And23660_o0 : std_logic;
	signal And23680_o0 : std_logic;
	signal And23700_o0 : std_logic;
	signal And23720_o0 : std_logic;
	signal And23740_o0 : std_logic;
	signal And23760_o0 : std_logic;
	signal And23780_o0 : std_logic;
	signal Or23800_o0 : std_logic;
	signal And23820_o0 : std_logic;
	signal Not3840_o0 : std_logic;
	signal Nand23860_o0 : std_logic;
	signal Or23880_o0 : std_logic;
	signal And23900_o0 : std_logic;
	signal And23920_o0 : std_logic;
	signal Or23940_o0 : std_logic;
	signal And23960_o0 : std_logic;
	signal Or23980_o0 : std_logic;
	signal Nor24000_o0 : std_logic;
	signal And24020_o0 : std_logic;
	signal And24040_o0 : std_logic;
	signal And24060_o0 : std_logic;
	signal And24080_o0 : std_logic;
	signal Or24100_o0 : std_logic;
	signal And24120_o0 : std_logic;
	signal And24140_o0 : std_logic;
	signal And24160_o0 : std_logic;
	signal And24180_o0 : std_logic;
	signal And24200_o0 : std_logic;
	signal And24220_o0 : std_logic;
	signal Or24240_o0 : std_logic;
	signal And24260_o0 : std_logic;
	signal And24280_o0 : std_logic;
	signal Nor24300_o0 : std_logic;
	signal And24320_o0 : std_logic;
	signal And24340_o0 : std_logic;
	signal Or24360_o0 : std_logic;
	signal And24380_o0 : std_logic;
	signal And24400_o0 : std_logic;
	signal And24420_o0 : std_logic;
	signal Or24440_o0 : std_logic;
	signal And24460_o0 : std_logic;
	signal And24480_o0 : std_logic;
	signal And24500_o0 : std_logic;
	signal Or24520_o0 : std_logic;
	signal And24540_o0 : std_logic;
	signal And24560_o0 : std_logic;
	signal And24580_o0 : std_logic;
	signal Or24600_o0 : std_logic;
	signal And24620_o0 : std_logic;
	signal And24640_o0 : std_logic;
	signal And24660_o0 : std_logic;
	signal Or24680_o0 : std_logic;
	signal And24700_o0 : std_logic;
	signal Or24720_o0 : std_logic;
	signal And24740_o0 : std_logic;
	signal And24760_o0 : std_logic;
	signal And24780_o0 : std_logic;
	signal And24800_o0 : std_logic;
	signal Or24820_o0 : std_logic;
	signal And24840_o0 : std_logic;
	signal And24860_o0 : std_logic;
	signal And24880_o0 : std_logic;
	signal And24900_o0 : std_logic;
	signal Nor24920_o0 : std_logic;
	signal And24940_o0 : std_logic;
	signal And24960_o0 : std_logic;
	signal And24980_o0 : std_logic;
	signal And25000_o0 : std_logic;
	signal And25020_o0 : std_logic;
	signal And25040_o0 : std_logic;
	signal Or25060_o0 : std_logic;
	signal And25080_o0 : std_logic;
	signal Nor25100_o0 : std_logic;
	signal And25120_o0 : std_logic;
	signal And25140_o0 : std_logic;
	signal Or25160_o0 : std_logic;
	signal And25180_o0 : std_logic;
	signal Xor25200_o0 : std_logic;
	signal Xor25220_o0 : std_logic;
	signal Nor25240_o0 : std_logic;
	signal And25260_o0 : std_logic;
	signal And25280_o0 : std_logic;
	signal And25300_o0 : std_logic;
	signal And25320_o0 : std_logic;
	signal And25340_o0 : std_logic;
	signal Or25360_o0 : std_logic;
	signal And25380_o0 : std_logic;
	signal Or25400_o0 : std_logic;
	signal And25420_o0 : std_logic;
	signal And25440_o0 : std_logic;
	signal And25460_o0 : std_logic;
	signal Or25480_o0 : std_logic;
	signal Or25500_o0 : std_logic;
	signal And25520_o0 : std_logic;
	signal Or25540_o0 : std_logic;
	signal Or25560_o0 : std_logic;
	signal And25580_o0 : std_logic;
	signal And25600_o0 : std_logic;
	signal And25620_o0 : std_logic;
	signal And25640_o0 : std_logic;
	signal Or25660_o0 : std_logic;
	signal And25680_o0 : std_logic;
	signal And25700_o0 : std_logic;
	signal And25720_o0 : std_logic;
	signal And25740_o0 : std_logic;
	signal And25760_o0 : std_logic;
	signal And25780_o0 : std_logic;
	signal And25800_o0 : std_logic;
	signal Or25820_o0 : std_logic;
	signal And25840_o0 : std_logic;
	signal And25860_o0 : std_logic;
	signal And25880_o0 : std_logic;
	signal Or25900_o0 : std_logic;
	signal And25920_o0 : std_logic;
	signal And25940_o0 : std_logic;
	signal And25960_o0 : std_logic;
	signal And25980_o0 : std_logic;
	signal Or26000_o0 : std_logic;
	signal And26020_o0 : std_logic;
	signal And26040_o0 : std_logic;
	signal And26060_o0 : std_logic;
	signal Or26080_o0 : std_logic;
	signal Or26100_o0 : std_logic;
	signal And26120_o0 : std_logic;
	signal And26140_o0 : std_logic;
	signal And26160_o0 : std_logic;
	signal And26180_o0 : std_logic;
	signal Or26200_o0 : std_logic;
	signal And26220_o0 : std_logic;
	signal And26240_o0 : std_logic;
	signal Or26260_o0 : std_logic;
	signal And26280_o0 : std_logic;
	signal And26300_o0 : std_logic;
	signal And26320_o0 : std_logic;
	signal Or26340_o0 : std_logic;
	signal And26360_o0 : std_logic;
	signal Or26380_o0 : std_logic;
	signal And26400_o0 : std_logic;
	signal And26420_o0 : std_logic;
	signal And26440_o0 : std_logic;
	signal And26460_o0 : std_logic;
	signal Or26480_o0 : std_logic;
	signal And26500_o0 : std_logic;
	signal And26520_o0 : std_logic;
	signal Xor26540_o0 : std_logic;
	signal Nor26560_o0 : std_logic;
	signal And26580_o0 : std_logic;
	signal And26600_o0 : std_logic;
	signal Or26620_o0 : std_logic;
	signal And26640_o0 : std_logic;
	signal Nor26660_o0 : std_logic;
	signal And26680_o0 : std_logic;
	signal And26700_o0 : std_logic;
	signal Or26720_o0 : std_logic;
	signal And26740_o0 : std_logic;
	signal And26760_o0 : std_logic;
	signal And26780_o0 : std_logic;
	signal And26800_o0 : std_logic;
	signal Or26820_o0 : std_logic;
	signal And26840_o0 : std_logic;
	signal And26860_o0 : std_logic;
	signal And26880_o0 : std_logic;
	signal And26900_o0 : std_logic;
	signal And26920_o0 : std_logic;
	signal Or26940_o0 : std_logic;
	signal And26960_o0 : std_logic;
	signal Xor26980_o0 : std_logic;
	signal Not7000_o0 : std_logic;
	signal And27020_o0 : std_logic;
	signal And27040_o0 : std_logic;
	signal And27060_o0 : std_logic;
	signal Or27080_o0 : std_logic;
	signal And27100_o0 : std_logic;
	signal Not7120_o0 : std_logic;
	signal Not7140_o0 : std_logic;
	signal Or27160_o0 : std_logic;
	signal Or27180_o0 : std_logic;
	signal Or27200_o0 : std_logic;
	signal And27220_o0 : std_logic;
	signal Or27240_o0 : std_logic;
	signal And27260_o0 : std_logic;
	signal Or27280_o0 : std_logic;
	signal And27300_o0 : std_logic;
	signal Or27320_o0 : std_logic;
	signal And27340_o0 : std_logic;
	signal Or27360_o0 : std_logic;
	signal And27380_o0 : std_logic;
	signal And27400_o0 : std_logic;
	signal And27420_o0 : std_logic;
	signal Not7440_o0 : std_logic;
	signal And27460_o0 : std_logic;
	signal Or27480_o0 : std_logic;
	signal And27500_o0 : std_logic;
	signal And27520_o0 : std_logic;
	signal And27540_o0 : std_logic;
	signal And27560_o0 : std_logic;
	signal Or27580_o0 : std_logic;
	signal Or27600_o0 : std_logic;
	signal And27620_o0 : std_logic;
	signal Or27640_o0 : std_logic;
	signal And27660_o0 : std_logic;
	signal And27680_o0 : std_logic;
	signal And27700_o0 : std_logic;
	signal Or27720_o0 : std_logic;
	signal And27740_o0 : std_logic;
	signal Or27760_o0 : std_logic;
	signal And27780_o0 : std_logic;
	signal Or27800_o0 : std_logic;
	signal And27820_o0 : std_logic;
	signal Nor27840_o0 : std_logic;
	signal And27860_o0 : std_logic;
	signal And27880_o0 : std_logic;
	signal Or27900_o0 : std_logic;
	signal And27920_o0 : std_logic;
	signal And27940_o0 : std_logic;
	signal And27960_o0 : std_logic;
	signal And27980_o0 : std_logic;
	signal Or28000_o0 : std_logic;
	signal And28020_o0 : std_logic;
	signal And28040_o0 : std_logic;
	signal And28060_o0 : std_logic;
	signal And28080_o0 : std_logic;
	signal And28100_o0 : std_logic;
	signal And28120_o0 : std_logic;
	signal And28140_o0 : std_logic;
	signal And28160_o0 : std_logic;
	signal And28180_o0 : std_logic;
	signal And28200_o0 : std_logic;
	signal Or28220_o0 : std_logic;
	signal And28240_o0 : std_logic;
	signal And28260_o0 : std_logic;
	signal And28280_o0 : std_logic;
	signal Or28300_o0 : std_logic;
	signal And28320_o0 : std_logic;
	signal And28340_o0 : std_logic;
	signal And28360_o0 : std_logic;
	signal Or28380_o0 : std_logic;
	signal And28400_o0 : std_logic;
	signal Or28420_o0 : std_logic;
	signal And28440_o0 : std_logic;
	signal And28460_o0 : std_logic;
	signal And28480_o0 : std_logic;
	signal And28500_o0 : std_logic;
	signal Or28520_o0 : std_logic;
	signal And28540_o0 : std_logic;
	signal And28560_o0 : std_logic;
	signal Or28580_o0 : std_logic;
	signal And28600_o0 : std_logic;
	signal And28620_o0 : std_logic;
	signal And28640_o0 : std_logic;
	signal Or28660_o0 : std_logic;
	signal And28680_o0 : std_logic;
	signal Or28700_o0 : std_logic;
	signal And28720_o0 : std_logic;
	signal Or28740_o0 : std_logic;
	signal And28760_o0 : std_logic;
	signal Or28780_o0 : std_logic;
	signal And28800_o0 : std_logic;
	signal Or28820_o0 : std_logic;
	signal And28840_o0 : std_logic;
	signal And28860_o0 : std_logic;
	signal And28880_o0 : std_logic;
	signal And28900_o0 : std_logic;
	signal And28920_o0 : std_logic;
	signal Or28940_o0 : std_logic;
	signal And28960_o0 : std_logic;
	signal And28980_o0 : std_logic;
	signal And29000_o0 : std_logic;
	signal Or29020_o0 : std_logic;
	signal And29040_o0 : std_logic;
	signal And29060_o0 : std_logic;
	signal And29080_o0 : std_logic;
	signal And29100_o0 : std_logic;
	signal Or29120_o0 : std_logic;
	signal And29140_o0 : std_logic;
	signal And29160_o0 : std_logic;
	signal And29180_o0 : std_logic;
	signal And29200_o0 : std_logic;
	signal And29220_o0 : std_logic;
	signal Or29240_o0 : std_logic;
	signal Nor29260_o0 : std_logic;
	signal And29280_o0 : std_logic;
	signal And29300_o0 : std_logic;
	signal And29320_o0 : std_logic;
	signal And29340_o0 : std_logic;
	signal And29360_o0 : std_logic;
	signal Or29380_o0 : std_logic;
	signal And29400_o0 : std_logic;
	signal And29420_o0 : std_logic;
	signal And29440_o0 : std_logic;
	signal Nor29460_o0 : std_logic;
	signal Or29480_o0 : std_logic;
	signal And29500_o0 : std_logic;
	signal And29520_o0 : std_logic;
	signal Not9540_o0 : std_logic;
	signal And29560_o0 : std_logic;
	signal Not9580_o0 : std_logic;
	signal Or29600_o0 : std_logic;
	signal And29620_o0 : std_logic;
	signal Nor29640_o0 : std_logic;
	signal Or29660_o0 : std_logic;
	signal And29680_o0 : std_logic;
	signal Not9700_o0 : std_logic;
	signal And29720_o0 : std_logic;
	signal And29740_o0 : std_logic;
	signal Or29760_o0 : std_logic;
	signal And29780_o0 : std_logic;
	signal Not9800_o0 : std_logic;
	signal And29820_o0 : std_logic;
	signal Or29840_o0 : std_logic;
	signal And29860_o0 : std_logic;
	signal And29880_o0 : std_logic;
	signal Or29900_o0 : std_logic;
	signal And29920_o0 : std_logic;
	signal And29940_o0 : std_logic;
	signal And29960_o0 : std_logic;
	signal Or29980_o0 : std_logic;
	signal And210000_o0 : std_logic;
	signal Nand210020_o0 : std_logic;
	signal And210040_o0 : std_logic;
	signal And210060_o0 : std_logic;
	signal Or210080_o0 : std_logic;
	signal And210100_o0 : std_logic;
	signal And210120_o0 : std_logic;
	signal Or210140_o0 : std_logic;
	signal And210160_o0 : std_logic;
	signal Or210180_o0 : std_logic;
	signal And210200_o0 : std_logic;
	signal Xor210220_o0 : std_logic;
	signal And210240_o0 : std_logic;
	signal And210260_o0 : std_logic;
	signal And210280_o0 : std_logic;
	signal Or210300_o0 : std_logic;
	signal Or210320_o0 : std_logic;
	signal And210340_o0 : std_logic;
	signal Or210360_o0 : std_logic;
	signal And210380_o0 : std_logic;
	signal Or210400_o0 : std_logic;
	signal And210420_o0 : std_logic;
	signal And210440_o0 : std_logic;
	signal Or210460_o0 : std_logic;
	signal And210480_o0 : std_logic;
	signal And210500_o0 : std_logic;
	signal Not10520_o0 : std_logic;
	signal And210540_o0 : std_logic;
	signal Nand210560_o0 : std_logic;
	signal And210580_o0 : std_logic;
	signal And210600_o0 : std_logic;
	signal Or210620_o0 : std_logic;
	signal Nand210640_o0 : std_logic;
	signal And210660_o0 : std_logic;
	signal And210680_o0 : std_logic;
	signal Or210700_o0 : std_logic;
	signal And210720_o0 : std_logic;
	signal And210740_o0 : std_logic;
	signal Or210760_o0 : std_logic;
	signal And210780_o0 : std_logic;
	signal And210800_o0 : std_logic;
	signal Or210820_o0 : std_logic;
	signal And210840_o0 : std_logic;
	signal And210860_o0 : std_logic;
	signal And210880_o0 : std_logic;
	signal Or210900_o0 : std_logic;
	signal And210920_o0 : std_logic;
	signal And210940_o0 : std_logic;
	signal And210960_o0 : std_logic;
	signal Or210980_o0 : std_logic;
	signal And211000_o0 : std_logic;
	signal And211020_o0 : std_logic;
	signal Nor211040_o0 : std_logic;
	signal And211060_o0 : std_logic;
	signal And211080_o0 : std_logic;
	signal Or211100_o0 : std_logic;
	signal Or211120_o0 : std_logic;
	signal And211140_o0 : std_logic;
	signal And211160_o0 : std_logic;
	signal And211180_o0 : std_logic;
	signal And211200_o0 : std_logic;
	signal And211220_o0 : std_logic;
	signal And211240_o0 : std_logic;
	signal And211260_o0 : std_logic;
	signal Or211280_o0 : std_logic;
	signal And211300_o0 : std_logic;
	signal Or211320_o0 : std_logic;
	signal And211340_o0 : std_logic;
	signal And211360_o0 : std_logic;
	signal Or211380_o0 : std_logic;
	signal And211400_o0 : std_logic;
	signal Or211420_o0 : std_logic;
	signal And211440_o0 : std_logic;
	signal And211460_o0 : std_logic;
	signal And211480_o0 : std_logic;
	signal Or211500_o0 : std_logic;
	signal And211520_o0 : std_logic;
	signal And211540_o0 : std_logic;
	signal Or211560_o0 : std_logic;
	signal And211580_o0 : std_logic;
	signal And211600_o0 : std_logic;
	signal And211620_o0 : std_logic;
	signal Or211640_o0 : std_logic;
	signal And211660_o0 : std_logic;
	signal And211680_o0 : std_logic;
	signal And211700_o0 : std_logic;
	signal Or211720_o0 : std_logic;
	signal And211740_o0 : std_logic;
	signal And211760_o0 : std_logic;
	signal Or211780_o0 : std_logic;
	signal And211800_o0 : std_logic;
	signal And211820_o0 : std_logic;
	signal Or211840_o0 : std_logic;
	signal And211860_o0 : std_logic;
	signal And211880_o0 : std_logic;
	signal Or211900_o0 : std_logic;
	signal And211920_o0 : std_logic;
	signal And211940_o0 : std_logic;
	signal And211960_o0 : std_logic;
	signal Or211980_o0 : std_logic;
	signal And212000_o0 : std_logic;
	signal And212020_o0 : std_logic;
	signal And212040_o0 : std_logic;
	signal Or212060_o0 : std_logic;
	signal And212080_o0 : std_logic;
	signal Not12100_o0 : std_logic;
	signal Not12120_o0 : std_logic;
	signal Or212140_o0 : std_logic;
	signal And212160_o0 : std_logic;
	signal And212180_o0 : std_logic;
	signal And212200_o0 : std_logic;
	signal And212220_o0 : std_logic;
	signal Not12240_o0 : std_logic;
	signal Nor212260_o0 : std_logic;
	signal And212280_o0 : std_logic;
	signal And212300_o0 : std_logic;
	signal Or212320_o0 : std_logic;
	signal And212340_o0 : std_logic;
	signal And212360_o0 : std_logic;
	signal And212380_o0 : std_logic;
	signal And212400_o0 : std_logic;
	signal And212420_o0 : std_logic;
	signal Or212440_o0 : std_logic;
	signal And212460_o0 : std_logic;
	signal And212480_o0 : std_logic;
	signal And212500_o0 : std_logic;
	signal Or212520_o0 : std_logic;
	signal And212540_o0 : std_logic;
	signal And212560_o0 : std_logic;
	signal And212580_o0 : std_logic;
	signal And212600_o0 : std_logic;
	signal Or212620_o0 : std_logic;
	signal Nor212640_o0 : std_logic;
	signal And212660_o0 : std_logic;
	signal And212680_o0 : std_logic;
	signal Nor212700_o0 : std_logic;
	signal And212720_o0 : std_logic;
	signal And212740_o0 : std_logic;
	signal And212760_o0 : std_logic;
	signal And212780_o0 : std_logic;
	signal Or212800_o0 : std_logic;
	signal And212820_o0 : std_logic;
	signal Not12840_o0 : std_logic;
	signal And212860_o0 : std_logic;
	signal And212880_o0 : std_logic;
	signal And212900_o0 : std_logic;
	signal And212920_o0 : std_logic;
	signal Nor212940_o0 : std_logic;
	signal Or212960_o0 : std_logic;
	signal And212980_o0 : std_logic;
	signal Or213000_o0 : std_logic;
	signal And213020_o0 : std_logic;
	signal And213040_o0 : std_logic;
	signal Or213060_o0 : std_logic;
	signal And213080_o0 : std_logic;
	signal And213100_o0 : std_logic;
	signal And213120_o0 : std_logic;
	signal Or213140_o0 : std_logic;
	signal And213160_o0 : std_logic;
	signal And213180_o0 : std_logic;
	signal And213200_o0 : std_logic;
	signal Or213220_o0 : std_logic;
	signal And213240_o0 : std_logic;
	signal And213260_o0 : std_logic;
	signal And213280_o0 : std_logic;
	signal And213300_o0 : std_logic;
	signal And213320_o0 : std_logic;
	signal Or213340_o0 : std_logic;
	signal And213360_o0 : std_logic;
	signal Nand213380_o0 : std_logic;
	signal Or213400_o0 : std_logic;
	signal And213420_o0 : std_logic;
	signal And213440_o0 : std_logic;
	signal Or213460_o0 : std_logic;
	signal And213480_o0 : std_logic;
	signal Or213500_o0 : std_logic;
	signal And213520_o0 : std_logic;
	signal And213540_o0 : std_logic;
	signal Or213560_o0 : std_logic;
	signal And213580_o0 : std_logic;
	signal And213600_o0 : std_logic;
	signal Or213620_o0 : std_logic;
	signal And213640_o0 : std_logic;
	signal Or213660_o0 : std_logic;
	signal And213680_o0 : std_logic;
	signal And213700_o0 : std_logic;
	signal And213720_o0 : std_logic;
	signal Or213740_o0 : std_logic;
	signal And213760_o0 : std_logic;
	signal Or213780_o0 : std_logic;
	signal And213800_o0 : std_logic;
	signal Not13820_o0 : std_logic;
	signal Nor213840_o0 : std_logic;
	signal Nand213860_o0 : std_logic;
	signal Or213880_o0 : std_logic;
	signal And213900_o0 : std_logic;
	signal And213920_o0 : std_logic;
	signal Or213940_o0 : std_logic;
	signal And213960_o0 : std_logic;
	signal And213980_o0 : std_logic;
	signal And214000_o0 : std_logic;
	signal Or214020_o0 : std_logic;
	signal And214040_o0 : std_logic;
	signal Or214060_o0 : std_logic;
	signal And214080_o0 : std_logic;
	signal And214100_o0 : std_logic;
	signal Nor214120_o0 : std_logic;
	signal And214140_o0 : std_logic;
	signal Or214160_o0 : std_logic;
	signal And214180_o0 : std_logic;
	signal And214200_o0 : std_logic;
	signal Or214220_o0 : std_logic;
	signal And214240_o0 : std_logic;
	signal And214260_o0 : std_logic;
	signal Or214280_o0 : std_logic;
	signal And214300_o0 : std_logic;
	signal And214320_o0 : std_logic;
	signal And214340_o0 : std_logic;
	signal And214360_o0 : std_logic;
	signal Or214380_o0 : std_logic;
	signal And214400_o0 : std_logic;
	signal And214420_o0 : std_logic;
	signal And214440_o0 : std_logic;
	signal And214460_o0 : std_logic;
	signal Or214480_o0 : std_logic;
	signal And214500_o0 : std_logic;
	signal And214520_o0 : std_logic;
	signal And214540_o0 : std_logic;
	signal And214560_o0 : std_logic;
	signal Or214580_o0 : std_logic;
	signal And214600_o0 : std_logic;
	signal And214620_o0 : std_logic;
	signal And214640_o0 : std_logic;
	signal And214660_o0 : std_logic;
	signal And214680_o0 : std_logic;
	signal And214700_o0 : std_logic;
	signal Or214720_o0 : std_logic;
	signal Nor214740_o0 : std_logic;
	signal And214760_o0 : std_logic;
	signal And214780_o0 : std_logic;
	signal And214800_o0 : std_logic;
	signal Or214820_o0 : std_logic;
	signal And214840_o0 : std_logic;
	signal And214860_o0 : std_logic;
	signal And214880_o0 : std_logic;
	signal Or214900_o0 : std_logic;
	signal And214920_o0 : std_logic;
	signal Or214940_o0 : std_logic;
	signal Nor214960_o0 : std_logic;
	signal Nor214980_o0 : std_logic;
	signal And215000_o0 : std_logic;
	signal And215020_o0 : std_logic;
	signal And215040_o0 : std_logic;
	signal And215060_o0 : std_logic;
	signal And215080_o0 : std_logic;
	signal And215100_o0 : std_logic;
	signal Or215120_o0 : std_logic;
	signal And215140_o0 : std_logic;
	signal And215160_o0 : std_logic;
	signal Or215180_o0 : std_logic;
	signal And215200_o0 : std_logic;
	signal And215220_o0 : std_logic;
	signal And215240_o0 : std_logic;
	signal Nor215260_o0 : std_logic;
	signal And215280_o0 : std_logic;
	signal And215300_o0 : std_logic;
	signal Or215320_o0 : std_logic;
	signal And215340_o0 : std_logic;
	signal And215360_o0 : std_logic;
	signal And215380_o0 : std_logic;
	signal Or215400_o0 : std_logic;
	signal And215420_o0 : std_logic;
	signal And215440_o0 : std_logic;
	signal And215460_o0 : std_logic;
	signal And215480_o0 : std_logic;
	signal Or215500_o0 : std_logic;
	signal And215520_o0 : std_logic;
	signal Or215540_o0 : std_logic;
	signal And215560_o0 : std_logic;
	signal And215580_o0 : std_logic;
	signal And215600_o0 : std_logic;
	signal Or215620_o0 : std_logic;
	signal And215640_o0 : std_logic;
	signal And215660_o0 : std_logic;
	signal Or215680_o0 : std_logic;
	signal Nor215700_o0 : std_logic;
	signal And215720_o0 : std_logic;
	signal And215740_o0 : std_logic;
	signal And215760_o0 : std_logic;
	signal Or215780_o0 : std_logic;
	signal And215800_o0 : std_logic;
	signal And215820_o0 : std_logic;
	signal And215840_o0 : std_logic;
	signal And215860_o0 : std_logic;
	signal Nor215880_o0 : std_logic;
	signal And215900_o0 : std_logic;
	signal Or215920_o0 : std_logic;
	signal And215940_o0 : std_logic;
	signal And215960_o0 : std_logic;
	signal And215980_o0 : std_logic;
	signal Or216000_o0 : std_logic;
	signal And216020_o0 : std_logic;
	signal And216040_o0 : std_logic;
	signal And216060_o0 : std_logic;
	signal And216080_o0 : std_logic;
	signal Or216100_o0 : std_logic;
	signal And216120_o0 : std_logic;
	signal Xor216140_o0 : std_logic;
	signal And216160_o0 : std_logic;
	signal Or216180_o0 : std_logic;
	signal And216200_o0 : std_logic;
	signal And216220_o0 : std_logic;
	signal Or216240_o0 : std_logic;
	signal And216260_o0 : std_logic;
	signal And216280_o0 : std_logic;
	signal And216300_o0 : std_logic;
	signal Or216320_o0 : std_logic;
	signal And216340_o0 : std_logic;
	signal Or216360_o0 : std_logic;
	signal And216380_o0 : std_logic;
	signal Nand216400_o0 : std_logic;
	signal And216420_o0 : std_logic;
	signal And216440_o0 : std_logic;
	signal Or216460_o0 : std_logic;
	signal And216480_o0 : std_logic;
	signal And216500_o0 : std_logic;
	signal And216520_o0 : std_logic;
	signal And216540_o0 : std_logic;
	signal And216560_o0 : std_logic;
	signal And216580_o0 : std_logic;
	signal And216600_o0 : std_logic;
	signal Or216620_o0 : std_logic;
	signal And216640_o0 : std_logic;
	signal And216660_o0 : std_logic;
	signal Or216680_o0 : std_logic;
	signal And216700_o0 : std_logic;
	signal And216720_o0 : std_logic;
	signal Or216740_o0 : std_logic;
	signal And216760_o0 : std_logic;
	signal Xor216780_o0 : std_logic;
	signal Not16800_o0 : std_logic;
	signal And216820_o0 : std_logic;
	signal Nand216840_o0 : std_logic;
	signal And216860_o0 : std_logic;
	signal Or216880_o0 : std_logic;
	signal And216900_o0 : std_logic;
	signal Or216920_o0 : std_logic;
	signal And216940_o0 : std_logic;
	signal And216960_o0 : std_logic;
	signal Or216980_o0 : std_logic;
	signal And217000_o0 : std_logic;
	signal Or217020_o0 : std_logic;
	signal And217040_o0 : std_logic;
	signal Or217060_o0 : std_logic;
	signal Or217080_o0 : std_logic;
	signal And217100_o0 : std_logic;
	signal And217120_o0 : std_logic;
	signal Or217140_o0 : std_logic;
	signal And217160_o0 : std_logic;
	signal And217180_o0 : std_logic;
	signal And217200_o0 : std_logic;
	signal Or217220_o0 : std_logic;
	signal And217240_o0 : std_logic;
	signal And217260_o0 : std_logic;
	signal And217280_o0 : std_logic;
	signal Or217300_o0 : std_logic;
	signal And217320_o0 : std_logic;
	signal And217340_o0 : std_logic;
	signal And217360_o0 : std_logic;
	signal Or217380_o0 : std_logic;
	signal And217400_o0 : std_logic;
	signal Nand217420_o0 : std_logic;
	signal And217440_o0 : std_logic;
	signal And217460_o0 : std_logic;
	signal Or217480_o0 : std_logic;
	signal And217500_o0 : std_logic;
	signal And217520_o0 : std_logic;
	signal Or217540_o0 : std_logic;
	signal Or217560_o0 : std_logic;
	signal And217580_o0 : std_logic;
	signal And217600_o0 : std_logic;
	signal Or217620_o0 : std_logic;
	signal And217640_o0 : std_logic;
	signal Or217660_o0 : std_logic;
	signal And217680_o0 : std_logic;
	signal And217700_o0 : std_logic;
	signal And217720_o0 : std_logic;
	signal Or217740_o0 : std_logic;
	signal And217760_o0 : std_logic;
	signal And217780_o0 : std_logic;
	signal And217800_o0 : std_logic;
	signal Or217820_o0 : std_logic;
	signal Xor217840_o0 : std_logic;
	signal And217860_o0 : std_logic;
	signal Nand217880_o0 : std_logic;
	signal Nor217900_o0 : std_logic;
	signal And217920_o0 : std_logic;
	signal And217940_o0 : std_logic;
	signal And217960_o0 : std_logic;
	signal Or217980_o0 : std_logic;
	signal And218000_o0 : std_logic;
	signal Xor218020_o0 : std_logic;
	signal Nor218040_o0 : std_logic;
	signal Or218060_o0 : std_logic;
	signal And218080_o0 : std_logic;
	signal And218100_o0 : std_logic;
	signal Or218120_o0 : std_logic;
	signal And218140_o0 : std_logic;
	signal And218160_o0 : std_logic;
	signal Or218180_o0 : std_logic;
	signal And218200_o0 : std_logic;
	signal Or218220_o0 : std_logic;
	signal And218240_o0 : std_logic;
	signal Nor218260_o0 : std_logic;
	signal And218280_o0 : std_logic;
	signal And218300_o0 : std_logic;
	signal Or218320_o0 : std_logic;
	signal And218340_o0 : std_logic;
	signal And218360_o0 : std_logic;
	signal Or218380_o0 : std_logic;
	signal And218400_o0 : std_logic;
	signal And218420_o0 : std_logic;
	signal And218440_o0 : std_logic;
	signal And218460_o0 : std_logic;
	signal And218480_o0 : std_logic;
	signal Or218500_o0 : std_logic;
	signal And218520_o0 : std_logic;
	signal And218540_o0 : std_logic;
	signal And218560_o0 : std_logic;
	signal And218580_o0 : std_logic;
	signal And218600_o0 : std_logic;
	signal Or218620_o0 : std_logic;
	signal And218640_o0 : std_logic;
	signal And218660_o0 : std_logic;
	signal And218680_o0 : std_logic;
	signal Or218700_o0 : std_logic;
	signal And218720_o0 : std_logic;
	signal And218740_o0 : std_logic;
	signal And218760_o0 : std_logic;
	signal Or218780_o0 : std_logic;
	signal And218800_o0 : std_logic;
	signal And218820_o0 : std_logic;
	signal And218840_o0 : std_logic;
	signal Or218860_o0 : std_logic;
	signal And218880_o0 : std_logic;
	signal And218900_o0 : std_logic;
	signal And218920_o0 : std_logic;
	signal Or218940_o0 : std_logic;
	signal And218960_o0 : std_logic;
	signal And218980_o0 : std_logic;
	signal And219000_o0 : std_logic;
	signal And219020_o0 : std_logic;
	signal And219040_o0 : std_logic;
	signal And219060_o0 : std_logic;
	signal And219080_o0 : std_logic;
	signal And219100_o0 : std_logic;
	signal And219120_o0 : std_logic;
	signal Or219140_o0 : std_logic;
	signal And219160_o0 : std_logic;
	signal Or219180_o0 : std_logic;
	signal Or219200_o0 : std_logic;
	signal And219220_o0 : std_logic;
	signal Or219240_o0 : std_logic;
	signal And219260_o0 : std_logic;
	signal Or219280_o0 : std_logic;
	signal And219300_o0 : std_logic;
	signal Or219320_o0 : std_logic;
	signal And219340_o0 : std_logic;
	signal Or219360_o0 : std_logic;
	signal And219380_o0 : std_logic;
	signal Or219400_o0 : std_logic;
	signal And219420_o0 : std_logic;
	signal And219440_o0 : std_logic;
	signal Or219460_o0 : std_logic;
	signal Or219480_o0 : std_logic;
	signal And219500_o0 : std_logic;
	signal And219520_o0 : std_logic;
	signal And219540_o0 : std_logic;
	signal Or219560_o0 : std_logic;
	signal And219580_o0 : std_logic;
	signal And219600_o0 : std_logic;
	signal And219620_o0 : std_logic;
	signal And219640_o0 : std_logic;
	signal Or219660_o0 : std_logic;
	signal And219680_o0 : std_logic;
	signal And219700_o0 : std_logic;
	signal Or219720_o0 : std_logic;
	signal And219740_o0 : std_logic;
	signal And219760_o0 : std_logic;
	signal And219780_o0 : std_logic;
	signal And219800_o0 : std_logic;
	signal And219820_o0 : std_logic;
	signal Or219840_o0 : std_logic;
	signal Or219860_o0 : std_logic;
	signal And219880_o0 : std_logic;
	signal And219900_o0 : std_logic;
	signal And219920_o0 : std_logic;
	signal And219940_o0 : std_logic;
	signal And219960_o0 : std_logic;
	signal And219980_o0 : std_logic;
	signal Or220000_o0 : std_logic;
	signal And220020_o0 : std_logic;
	signal And220040_o0 : std_logic;
	signal Nor220060_o0 : std_logic;
	signal And220080_o0 : std_logic;
	signal And220100_o0 : std_logic;
	signal And220120_o0 : std_logic;
	signal Or220140_o0 : std_logic;
	signal And220160_o0 : std_logic;
	signal And220180_o0 : std_logic;
	signal And220200_o0 : std_logic;
	signal And220220_o0 : std_logic;
	signal And220240_o0 : std_logic;
	signal Or220260_o0 : std_logic;
	signal And220280_o0 : std_logic;
	signal Or220300_o0 : std_logic;
	signal Or220320_o0 : std_logic;
	signal Nor220340_o0 : std_logic;
	signal And220360_o0 : std_logic;
	signal And220380_o0 : std_logic;
	signal And220400_o0 : std_logic;
	signal And220420_o0 : std_logic;
	signal And220440_o0 : std_logic;
	signal And220460_o0 : std_logic;
	signal Or220480_o0 : std_logic;
	signal And220500_o0 : std_logic;
	signal Not20520_o0 : std_logic;
	signal And220540_o0 : std_logic;
	signal And220560_o0 : std_logic;
	signal And220580_o0 : std_logic;
	signal And220600_o0 : std_logic;
	signal Or220620_o0 : std_logic;
	signal And220640_o0 : std_logic;
	signal And220660_o0 : std_logic;
	signal And220680_o0 : std_logic;
	signal Or220700_o0 : std_logic;
	signal Or220720_o0 : std_logic;
	signal And220740_o0 : std_logic;
	signal Not20760_o0 : std_logic;
	signal Or220780_o0 : std_logic;
	signal And220800_o0 : std_logic;
	signal And220820_o0 : std_logic;
	signal Or220840_o0 : std_logic;
	signal And220860_o0 : std_logic;
	signal Or220880_o0 : std_logic;
	signal And220900_o0 : std_logic;
	signal Or220920_o0 : std_logic;
	signal And220940_o0 : std_logic;
	signal And220960_o0 : std_logic;
	signal Or220980_o0 : std_logic;
	signal And221000_o0 : std_logic;
	signal Xor221020_o0 : std_logic;
	signal Or221040_o0 : std_logic;
	signal And221060_o0 : std_logic;
	signal And221080_o0 : std_logic;
	signal Or221100_o0 : std_logic;
	signal And221120_o0 : std_logic;
	signal And221140_o0 : std_logic;
	signal Or221160_o0 : std_logic;
	signal And221180_o0 : std_logic;
	signal Or221200_o0 : std_logic;
	signal And221220_o0 : std_logic;
	signal And221240_o0 : std_logic;
	signal Or221260_o0 : std_logic;
	signal And221280_o0 : std_logic;
	signal Or221300_o0 : std_logic;
	signal And221320_o0 : std_logic;
	signal Nand221340_o0 : std_logic;
	signal And221360_o0 : std_logic;
	signal And221380_o0 : std_logic;
	signal Or221400_o0 : std_logic;
	signal And221420_o0 : std_logic;
	signal And221440_o0 : std_logic;
	signal And221460_o0 : std_logic;
	signal And221480_o0 : std_logic;
	signal Or221500_o0 : std_logic;
	signal And221520_o0 : std_logic;
	signal Or221540_o0 : std_logic;
	signal And221560_o0 : std_logic;
	signal Or221580_o0 : std_logic;
	signal And221600_o0 : std_logic;
	signal And221620_o0 : std_logic;
	signal And221640_o0 : std_logic;
	signal Or221660_o0 : std_logic;
	signal And221680_o0 : std_logic;
	signal And221700_o0 : std_logic;
	signal And221720_o0 : std_logic;
	signal And221740_o0 : std_logic;
	signal Or221760_o0 : std_logic;
	signal And221780_o0 : std_logic;
	signal And221800_o0 : std_logic;
	signal Or221820_o0 : std_logic;
	signal And221840_o0 : std_logic;
	signal And221860_o0 : std_logic;
	signal And221880_o0 : std_logic;
	signal Or221900_o0 : std_logic;
	signal Nor221920_o0 : std_logic;
	signal And221940_o0 : std_logic;
	signal And221960_o0 : std_logic;
	signal Or221980_o0 : std_logic;
	signal And222000_o0 : std_logic;
	signal And222020_o0 : std_logic;
	signal And222040_o0 : std_logic;
	signal Or222060_o0 : std_logic;
	signal And222080_o0 : std_logic;
	signal And222100_o0 : std_logic;
	signal And222120_o0 : std_logic;
	signal And222140_o0 : std_logic;
	signal And222160_o0 : std_logic;
	signal And222180_o0 : std_logic;
	signal Or222200_o0 : std_logic;
	signal And222220_o0 : std_logic;
	signal And222240_o0 : std_logic;
	signal And222260_o0 : std_logic;
	signal Or222280_o0 : std_logic;
	signal And222300_o0 : std_logic;
	signal And222320_o0 : std_logic;
	signal And222340_o0 : std_logic;
	signal Or222360_o0 : std_logic;
	signal And222380_o0 : std_logic;
	signal And222400_o0 : std_logic;
	signal Or222420_o0 : std_logic;
	signal And222440_o0 : std_logic;
	signal And222460_o0 : std_logic;
	signal And222480_o0 : std_logic;
	signal And222500_o0 : std_logic;
	signal And222520_o0 : std_logic;
	signal And222540_o0 : std_logic;
	signal Or222560_o0 : std_logic;
	signal Or222580_o0 : std_logic;
	signal Or222600_o0 : std_logic;
	signal And222620_o0 : std_logic;
	signal Or222640_o0 : std_logic;
	signal And222660_o0 : std_logic;
	signal And222680_o0 : std_logic;
	signal And222700_o0 : std_logic;
	signal And222720_o0 : std_logic;
	signal Or222740_o0 : std_logic;
	signal And222760_o0 : std_logic;
	signal And222780_o0 : std_logic;
	signal And222800_o0 : std_logic;
	signal And222820_o0 : std_logic;
	signal And222840_o0 : std_logic;
	signal And222860_o0 : std_logic;
	signal Nor222880_o0 : std_logic;
	signal And222900_o0 : std_logic;
	signal And222920_o0 : std_logic;
	signal And222940_o0 : std_logic;
	signal Or222960_o0 : std_logic;
	signal And222980_o0 : std_logic;
	signal Or223000_o0 : std_logic;
	signal And223020_o0 : std_logic;
	signal Or223040_o0 : std_logic;
	signal And223060_o0 : std_logic;
	signal And223080_o0 : std_logic;
	signal And223100_o0 : std_logic;
	signal Or223120_o0 : std_logic;
	signal And223140_o0 : std_logic;
	signal And223160_o0 : std_logic;
	signal And223180_o0 : std_logic;
	signal Or223200_o0 : std_logic;
	signal And223220_o0 : std_logic;
	signal And223240_o0 : std_logic;
	signal And223260_o0 : std_logic;
	signal And223280_o0 : std_logic;
	signal And223300_o0 : std_logic;
	signal Or223320_o0 : std_logic;
	signal And223340_o0 : std_logic;
	signal Or223360_o0 : std_logic;
	signal And223380_o0 : std_logic;
	signal And223400_o0 : std_logic;
	signal And223420_o0 : std_logic;
	signal And223440_o0 : std_logic;
	signal Or223460_o0 : std_logic;
	signal And223480_o0 : std_logic;
	signal And223500_o0 : std_logic;
	signal And223520_o0 : std_logic;
	signal And223540_o0 : std_logic;
	signal Or223560_o0 : std_logic;
	signal And223580_o0 : std_logic;
	signal And223600_o0 : std_logic;
	signal And223620_o0 : std_logic;
	signal And223640_o0 : std_logic;
	signal Or223660_o0 : std_logic;
	signal And223680_o0 : std_logic;
	signal And223700_o0 : std_logic;
	signal Or223720_o0 : std_logic;
	signal And223740_o0 : std_logic;
	signal And223760_o0 : std_logic;
	signal Nand223780_o0 : std_logic;
	signal And223800_o0 : std_logic;
	signal And223820_o0 : std_logic;
	signal Or223840_o0 : std_logic;
	signal And223860_o0 : std_logic;
	signal And223880_o0 : std_logic;
	signal And223900_o0 : std_logic;
	signal Or223920_o0 : std_logic;
	signal And223940_o0 : std_logic;
	signal Or223960_o0 : std_logic;
	signal And223980_o0 : std_logic;
	signal Nor224000_o0 : std_logic;
	signal And224020_o0 : std_logic;
	signal Or224040_o0 : std_logic;
	signal And224060_o0 : std_logic;
	signal And224080_o0 : std_logic;
	signal And224100_o0 : std_logic;
	signal Or224120_o0 : std_logic;
	signal And224140_o0 : std_logic;
	signal And224160_o0 : std_logic;
	signal And224180_o0 : std_logic;
	signal And224200_o0 : std_logic;
	signal And224220_o0 : std_logic;
	signal And224240_o0 : std_logic;
	signal And224260_o0 : std_logic;
	signal Or224280_o0 : std_logic;
	signal And224300_o0 : std_logic;
	signal And224320_o0 : std_logic;
	signal And224340_o0 : std_logic;
	signal And224360_o0 : std_logic;
	signal And224380_o0 : std_logic;
	signal And224400_o0 : std_logic;
	signal Or224420_o0 : std_logic;
	signal And224440_o0 : std_logic;
	signal And224460_o0 : std_logic;
	signal And224480_o0 : std_logic;
	signal And224500_o0 : std_logic;
	signal And224520_o0 : std_logic;
	signal And224540_o0 : std_logic;
	signal Not24560_o0 : std_logic;
	signal And224580_o0 : std_logic;
	signal And224600_o0 : std_logic;
	signal And224620_o0 : std_logic;
	signal And224640_o0 : std_logic;
	signal And224660_o0 : std_logic;
	signal Or224680_o0 : std_logic;
	signal And224700_o0 : std_logic;
	signal And224720_o0 : std_logic;
	signal And224740_o0 : std_logic;
	signal Or224760_o0 : std_logic;
	signal Or224780_o0 : std_logic;
	signal Or224800_o0 : std_logic;
	signal Or224820_o0 : std_logic;
	signal And224840_o0 : std_logic;
	signal Or224860_o0 : std_logic;
	signal And224880_o0 : std_logic;
	signal And224900_o0 : std_logic;
	signal Or224920_o0 : std_logic;
	signal Or224940_o0 : std_logic;
	signal Not24960_o0 : std_logic;
	signal And224980_o0 : std_logic;
	signal And225000_o0 : std_logic;
	signal Or225020_o0 : std_logic;
	signal And225040_o0 : std_logic;
	signal And225060_o0 : std_logic;
	signal And225080_o0 : std_logic;
	signal Or225100_o0 : std_logic;
	signal And225120_o0 : std_logic;
	signal And225140_o0 : std_logic;
	signal And225160_o0 : std_logic;
	signal Or225180_o0 : std_logic;
	signal And225200_o0 : std_logic;
	signal And225220_o0 : std_logic;
	signal And225240_o0 : std_logic;
	signal And225260_o0 : std_logic;
	signal Or225280_o0 : std_logic;
	signal And225300_o0 : std_logic;
	signal And225320_o0 : std_logic;
	signal And225340_o0 : std_logic;
	signal Or225360_o0 : std_logic;
	signal And225380_o0 : std_logic;
	signal And225400_o0 : std_logic;
	signal Or225420_o0 : std_logic;
	signal And225440_o0 : std_logic;
	signal And225460_o0 : std_logic;
	signal Or225480_o0 : std_logic;
	signal And225500_o0 : std_logic;
	signal And225520_o0 : std_logic;
	signal Or225540_o0 : std_logic;
	signal And225560_o0 : std_logic;
	signal And225580_o0 : std_logic;
	signal And225600_o0 : std_logic;
	signal And225620_o0 : std_logic;
	signal Or225640_o0 : std_logic;
	signal And225660_o0 : std_logic;
	signal And225680_o0 : std_logic;
	signal And225700_o0 : std_logic;
	signal And225720_o0 : std_logic;
	signal Or225740_o0 : std_logic;
	signal And225760_o0 : std_logic;
	signal And225780_o0 : std_logic;
	signal And225800_o0 : std_logic;
	signal And225820_o0 : std_logic;
	signal Or225840_o0 : std_logic;
	signal Nor225860_o0 : std_logic;
	signal And225880_o0 : std_logic;
	signal And225900_o0 : std_logic;
	signal And225920_o0 : std_logic;
	signal Or225940_o0 : std_logic;
	signal And225960_o0 : std_logic;
	signal And225980_o0 : std_logic;
	signal And226000_o0 : std_logic;
	signal Nor226020_o0 : std_logic;
	signal And226040_o0 : std_logic;
	signal And226060_o0 : std_logic;
	signal And226080_o0 : std_logic;
	signal And226100_o0 : std_logic;
	signal Or226120_o0 : std_logic;
	signal Nor226140_o0 : std_logic;
	signal Nor226160_o0 : std_logic;
	signal And226180_o0 : std_logic;
	signal And226200_o0 : std_logic;
	signal And226220_o0 : std_logic;
	signal Or226240_o0 : std_logic;
	signal And226260_o0 : std_logic;
	signal And226280_o0 : std_logic;
	signal Or226300_o0 : std_logic;
	signal And226320_o0 : std_logic;
	signal And226340_o0 : std_logic;
	signal And226360_o0 : std_logic;
	signal Or226380_o0 : std_logic;
	signal And226400_o0 : std_logic;
	signal And226420_o0 : std_logic;
	signal And226440_o0 : std_logic;
	signal Or226460_o0 : std_logic;
	signal And226480_o0 : std_logic;
	signal Nor226500_o0 : std_logic;
	signal And226520_o0 : std_logic;
	signal And226540_o0 : std_logic;
	signal And226560_o0 : std_logic;
	signal Or226580_o0 : std_logic;
	signal And226600_o0 : std_logic;
	signal And226620_o0 : std_logic;
	signal And226640_o0 : std_logic;
	signal Or226660_o0 : std_logic;
	signal And226680_o0 : std_logic;
	signal Or226700_o0 : std_logic;
	signal And226720_o0 : std_logic;
	signal Xor226740_o0 : std_logic;
	signal And226760_o0 : std_logic;
	signal And226780_o0 : std_logic;
	signal And226800_o0 : std_logic;
	signal Or226820_o0 : std_logic;
	signal And226840_o0 : std_logic;
	signal Or226860_o0 : std_logic;
	signal And226880_o0 : std_logic;
	signal Or226900_o0 : std_logic;
	signal And226920_o0 : std_logic;
	signal And226940_o0 : std_logic;
	signal And226960_o0 : std_logic;
	signal Or226980_o0 : std_logic;
	signal And227000_o0 : std_logic;
	signal And227020_o0 : std_logic;
	signal And227040_o0 : std_logic;
	signal And227060_o0 : std_logic;
	signal Or227080_o0 : std_logic;
	signal And227100_o0 : std_logic;
	signal And227120_o0 : std_logic;
	signal Or227140_o0 : std_logic;
	signal And227160_o0 : std_logic;
	signal And227180_o0 : std_logic;
	signal And227200_o0 : std_logic;
	signal And227220_o0 : std_logic;
	signal And227240_o0 : std_logic;
	signal And227260_o0 : std_logic;
	signal And227280_o0 : std_logic;
	signal And227300_o0 : std_logic;
	signal And227320_o0 : std_logic;
	signal Or227340_o0 : std_logic;
	signal Or227360_o0 : std_logic;
	signal Or227380_o0 : std_logic;
	signal And227400_o0 : std_logic;
	signal And227420_o0 : std_logic;
	signal And227440_o0 : std_logic;
	signal And227460_o0 : std_logic;
	signal Or227480_o0 : std_logic;
	signal And227500_o0 : std_logic;
	signal And227520_o0 : std_logic;
	signal And227540_o0 : std_logic;
	signal Or227560_o0 : std_logic;
	signal And227580_o0 : std_logic;
	signal And227600_o0 : std_logic;
	signal And227620_o0 : std_logic;
	signal And227640_o0 : std_logic;
	signal Or227660_o0 : std_logic;
	signal And227680_o0 : std_logic;
	signal Or227700_o0 : std_logic;
	signal Nor227720_o0 : std_logic;
	signal And227740_o0 : std_logic;
	signal Or227760_o0 : std_logic;
	signal And227780_o0 : std_logic;
	signal Xor227800_o0 : std_logic;
	signal Not27820_o0 : std_logic;
	signal And227840_o0 : std_logic;
	signal Or227860_o0 : std_logic;
	signal Or227880_o0 : std_logic;
	signal And227900_o0 : std_logic;
	signal Or227920_o0 : std_logic;
	signal And227940_o0 : std_logic;
	signal Or227960_o0 : std_logic;
	signal And227980_o0 : std_logic;
	signal Or228000_o0 : std_logic;
	signal And228020_o0 : std_logic;
	signal And228040_o0 : std_logic;
	signal Or228060_o0 : std_logic;
	signal And228080_o0 : std_logic;
	signal Or228100_o0 : std_logic;
	signal And228120_o0 : std_logic;
	signal Xor228140_o0 : std_logic;
	signal Not28160_o0 : std_logic;
	signal Or228180_o0 : std_logic;
	signal And228200_o0 : std_logic;
	signal Or228220_o0 : std_logic;
	signal And228240_o0 : std_logic;
	signal And228260_o0 : std_logic;
	signal And228280_o0 : std_logic;
	signal Or228300_o0 : std_logic;
	signal And228320_o0 : std_logic;
	signal And228340_o0 : std_logic;
	signal Or228360_o0 : std_logic;
	signal And228380_o0 : std_logic;
	signal Or228400_o0 : std_logic;
	signal And228420_o0 : std_logic;
	signal Or228440_o0 : std_logic;
	signal Or228460_o0 : std_logic;
	signal And228480_o0 : std_logic;
	signal Or228500_o0 : std_logic;
	signal And228520_o0 : std_logic;
	signal Or228540_o0 : std_logic;
	signal And228560_o0 : std_logic;
	signal And228580_o0 : std_logic;
	signal And228600_o0 : std_logic;
	signal Or228620_o0 : std_logic;
	signal And228640_o0 : std_logic;
	signal And228660_o0 : std_logic;
	signal And228680_o0 : std_logic;
	signal Or228700_o0 : std_logic;
	signal And228720_o0 : std_logic;
	signal And228740_o0 : std_logic;
	signal And228760_o0 : std_logic;
	signal Or228780_o0 : std_logic;
	signal Or228800_o0 : std_logic;
	signal And228820_o0 : std_logic;
	signal And228840_o0 : std_logic;
	signal Or228860_o0 : std_logic;
	signal And228880_o0 : std_logic;
	signal And228900_o0 : std_logic;
	signal Or228920_o0 : std_logic;
	signal And228940_o0 : std_logic;
	signal And228960_o0 : std_logic;
	signal And228980_o0 : std_logic;
	signal Or229000_o0 : std_logic;
	signal And229020_o0 : std_logic;
	signal And229040_o0 : std_logic;
	signal And229060_o0 : std_logic;
	signal Or229080_o0 : std_logic;
	signal And229100_o0 : std_logic;
	signal Or229120_o0 : std_logic;
	signal Or229140_o0 : std_logic;
	signal Or229160_o0 : std_logic;
	signal And229180_o0 : std_logic;
	signal Or229200_o0 : std_logic;
	signal And229220_o0 : std_logic;
	signal And229240_o0 : std_logic;
	signal Or229260_o0 : std_logic;
	signal Nor229280_o0 : std_logic;
	signal And229300_o0 : std_logic;
	signal And229320_o0 : std_logic;
	signal And229340_o0 : std_logic;
	signal And229360_o0 : std_logic;
	signal And229380_o0 : std_logic;
	signal Or229400_o0 : std_logic;
	signal And229420_o0 : std_logic;
	signal And229440_o0 : std_logic;
	signal Or229460_o0 : std_logic;
	signal And229480_o0 : std_logic;
	signal Nor229500_o0 : std_logic;
	signal Or229520_o0 : std_logic;
	signal And229540_o0 : std_logic;
	signal Or229560_o0 : std_logic;
	signal And229580_o0 : std_logic;
	signal And229600_o0 : std_logic;
	signal And229620_o0 : std_logic;
	signal Or229640_o0 : std_logic;
	signal And229660_o0 : std_logic;
	signal Or229680_o0 : std_logic;
	signal And229700_o0 : std_logic;
	signal And229720_o0 : std_logic;
	signal Or229740_o0 : std_logic;
	signal And229760_o0 : std_logic;
	signal Or229780_o0 : std_logic;
	signal And229800_o0 : std_logic;
	signal And229820_o0 : std_logic;
	signal Or229840_o0 : std_logic;
	signal And229860_o0 : std_logic;
	signal And229880_o0 : std_logic;
	signal Or229900_o0 : std_logic;
	signal And229920_o0 : std_logic;
	signal And229940_o0 : std_logic;
	signal Or229960_o0 : std_logic;
	signal And229980_o0 : std_logic;
	signal And230000_o0 : std_logic;
	signal Nor230020_o0 : std_logic;
	signal And230040_o0 : std_logic;
	signal Or230060_o0 : std_logic;
	signal And230080_o0 : std_logic;
	signal And230100_o0 : std_logic;
	signal Or230120_o0 : std_logic;
	signal And230140_o0 : std_logic;
	signal Or230160_o0 : std_logic;
	signal And230180_o0 : std_logic;
	signal And230200_o0 : std_logic;
	signal Or230220_o0 : std_logic;
	signal And230240_o0 : std_logic;
	signal And230260_o0 : std_logic;
	signal Or230280_o0 : std_logic;
	signal And230300_o0 : std_logic;
	signal And230320_o0 : std_logic;
	signal And230340_o0 : std_logic;
	signal And230360_o0 : std_logic;
	signal And230380_o0 : std_logic;
	signal And230400_o0 : std_logic;
	signal And230420_o0 : std_logic;
	signal Or230440_o0 : std_logic;
	signal And230460_o0 : std_logic;
	signal And230480_o0 : std_logic;
	signal And230500_o0 : std_logic;
	signal And230520_o0 : std_logic;
	signal And230540_o0 : std_logic;
	signal And230560_o0 : std_logic;
	signal And230580_o0 : std_logic;
	signal Or230600_o0 : std_logic;
	signal And230620_o0 : std_logic;
	signal And230640_o0 : std_logic;
	signal Or230660_o0 : std_logic;
	signal And230680_o0 : std_logic;
	signal And230700_o0 : std_logic;
	signal And230720_o0 : std_logic;
	signal And230740_o0 : std_logic;
	signal And230760_o0 : std_logic;
	signal And230780_o0 : std_logic;
	signal And230800_o0 : std_logic;
	signal Or230820_o0 : std_logic;
	signal Or230840_o0 : std_logic;
	signal And230860_o0 : std_logic;
	signal And230880_o0 : std_logic;
	signal Or230900_o0 : std_logic;
	signal And230920_o0 : std_logic;
	signal Or230940_o0 : std_logic;
	signal And230960_o0 : std_logic;
	signal And230980_o0 : std_logic;
	signal And231000_o0 : std_logic;
	signal Or231020_o0 : std_logic;
	signal And231040_o0 : std_logic;
	signal And231060_o0 : std_logic;
	signal And231080_o0 : std_logic;
	signal Or231100_o0 : std_logic;
	signal And231120_o0 : std_logic;
	signal And231140_o0 : std_logic;
	signal And231160_o0 : std_logic;
	signal Or231180_o0 : std_logic;
	signal And231200_o0 : std_logic;
	signal And231220_o0 : std_logic;
	signal And231240_o0 : std_logic;
	signal And231260_o0 : std_logic;
	signal Or231280_o0 : std_logic;
	signal Or231300_o0 : std_logic;
	signal And231320_o0 : std_logic;
	signal And231340_o0 : std_logic;
	signal And231360_o0 : std_logic;
	signal And231380_o0 : std_logic;
	signal And231400_o0 : std_logic;
	signal And231420_o0 : std_logic;
	signal And231440_o0 : std_logic;
	signal Or231460_o0 : std_logic;
	signal And231480_o0 : std_logic;
	signal Or231500_o0 : std_logic;
	signal And231520_o0 : std_logic;
	signal And231540_o0 : std_logic;
	signal Or231560_o0 : std_logic;
	signal And231580_o0 : std_logic;
	signal And231600_o0 : std_logic;
	signal Or231620_o0 : std_logic;
	signal And231640_o0 : std_logic;
	signal Or231660_o0 : std_logic;
	signal And231680_o0 : std_logic;
	signal Nand231700_o0 : std_logic;
	signal Or231720_o0 : std_logic;
	signal And231740_o0 : std_logic;
	signal Or231760_o0 : std_logic;
	signal And231780_o0 : std_logic;
	signal And231800_o0 : std_logic;
	signal Or231820_o0 : std_logic;
	signal And231840_o0 : std_logic;
	signal Or231860_o0 : std_logic;
	signal Or231880_o0 : std_logic;
	signal And231900_o0 : std_logic;
	signal And231920_o0 : std_logic;
	signal Or231940_o0 : std_logic;
	signal And231960_o0 : std_logic;
	signal Or231980_o0 : std_logic;
	signal And232000_o0 : std_logic;
	signal And232020_o0 : std_logic;
	signal Or232040_o0 : std_logic;
	signal And232060_o0 : std_logic;
	signal Nand232080_o0 : std_logic;
	signal And232100_o0 : std_logic;
	signal Or232120_o0 : std_logic;
	signal And232140_o0 : std_logic;
	signal And232160_o0 : std_logic;
	signal And232180_o0 : std_logic;
	signal And232200_o0 : std_logic;
	signal Nor232220_o0 : std_logic;
	signal And232240_o0 : std_logic;
	signal Or232260_o0 : std_logic;
	signal Or232280_o0 : std_logic;
	signal Or232300_o0 : std_logic;
	signal And232320_o0 : std_logic;
	signal Or232340_o0 : std_logic;
	signal And232360_o0 : std_logic;
	signal And232380_o0 : std_logic;
	signal And232400_o0 : std_logic;
	signal And232420_o0 : std_logic;
	signal And232440_o0 : std_logic;
	signal Or232460_o0 : std_logic;
	signal Or232480_o0 : std_logic;
	signal And232500_o0 : std_logic;
	signal And232520_o0 : std_logic;
	signal Or232540_o0 : std_logic;
	signal And232560_o0 : std_logic;
	signal Or232580_o0 : std_logic;
	signal And232600_o0 : std_logic;
	signal Not32620_o0 : std_logic;
	signal And232640_o0 : std_logic;
	signal And232660_o0 : std_logic;
	signal Or232680_o0 : std_logic;
	signal And232700_o0 : std_logic;
	signal Or232720_o0 : std_logic;
	signal And232740_o0 : std_logic;
	signal And232760_o0 : std_logic;
	signal Or232780_o0 : std_logic;
	signal Or232800_o0 : std_logic;
	signal And232820_o0 : std_logic;
	signal Or232840_o0 : std_logic;
	signal And232860_o0 : std_logic;
	signal And232880_o0 : std_logic;
	signal Or232900_o0 : std_logic;
	signal Or232920_o0 : std_logic;
	signal And232940_o0 : std_logic;
	signal Or232960_o0 : std_logic;
	signal And232980_o0 : std_logic;
	signal And233000_o0 : std_logic;
	signal Or233020_o0 : std_logic;
	signal And233040_o0 : std_logic;
	signal Or233060_o0 : std_logic;
	signal And233080_o0 : std_logic;
	signal And233100_o0 : std_logic;
	signal Or233120_o0 : std_logic;
	signal Or233140_o0 : std_logic;
	signal And233160_o0 : std_logic;
	signal And233180_o0 : std_logic;
	signal Or233200_o0 : std_logic;
	signal And233220_o0 : std_logic;
	signal And233240_o0 : std_logic;
	signal Or233260_o0 : std_logic;
	signal And233280_o0 : std_logic;
	signal Nor233300_o0 : std_logic;
	signal Or233320_o0 : std_logic;
	signal Or233340_o0 : std_logic;
	signal And233360_o0 : std_logic;
	signal And233380_o0 : std_logic;
	signal And233400_o0 : std_logic;
	signal Or233420_o0 : std_logic;
	signal And233440_o0 : std_logic;
	signal Or233460_o0 : std_logic;
	signal And233480_o0 : std_logic;
	signal And233500_o0 : std_logic;
	signal And233520_o0 : std_logic;
	signal And233540_o0 : std_logic;
	signal Or233560_o0 : std_logic;
	signal And233580_o0 : std_logic;
	signal And233600_o0 : std_logic;
	signal Or233620_o0 : std_logic;
	signal And233640_o0 : std_logic;
	signal And233660_o0 : std_logic;
	signal And233680_o0 : std_logic;
	signal Or233700_o0 : std_logic;
	signal And233720_o0 : std_logic;
	signal And233740_o0 : std_logic;
	signal And233760_o0 : std_logic;
	signal Or233780_o0 : std_logic;
	signal And233800_o0 : std_logic;
	signal Or233820_o0 : std_logic;
	signal Or233840_o0 : std_logic;
	signal Or233860_o0 : std_logic;
	signal And233880_o0 : std_logic;
	signal Or233900_o0 : std_logic;
	signal And233920_o0 : std_logic;
	signal And233940_o0 : std_logic;
	signal And233960_o0 : std_logic;
	signal Or233980_o0 : std_logic;
	signal And234000_o0 : std_logic;
	signal Or234020_o0 : std_logic;
	signal And234040_o0 : std_logic;
	signal And234060_o0 : std_logic;
	signal And234080_o0 : std_logic;
	signal Or234100_o0 : std_logic;
	signal And234120_o0 : std_logic;
	signal Nor234140_o0 : std_logic;
	signal And234160_o0 : std_logic;
	signal And234180_o0 : std_logic;
	signal And234200_o0 : std_logic;
	signal Or234220_o0 : std_logic;
	signal Or234240_o0 : std_logic;
	signal And234260_o0 : std_logic;
	signal And234280_o0 : std_logic;
	signal And234300_o0 : std_logic;
	signal And234320_o0 : std_logic;
	signal Or234340_o0 : std_logic;
	signal And234360_o0 : std_logic;
	signal And234380_o0 : std_logic;
	signal And234400_o0 : std_logic;
	signal And234420_o0 : std_logic;
	signal Or234440_o0 : std_logic;
	signal And234460_o0 : std_logic;
	signal And234480_o0 : std_logic;
	signal Or234500_o0 : std_logic;
	signal And234520_o0 : std_logic;
	signal And234540_o0 : std_logic;
	signal And234560_o0 : std_logic;
	signal And234580_o0 : std_logic;
	signal And234600_o0 : std_logic;
	signal And234620_o0 : std_logic;
	signal And234640_o0 : std_logic;
	signal And234660_o0 : std_logic;
	signal And234680_o0 : std_logic;
	signal Or234700_o0 : std_logic;
	signal And234720_o0 : std_logic;
	signal And234740_o0 : std_logic;
	signal And234760_o0 : std_logic;
	signal And234780_o0 : std_logic;
	signal And234800_o0 : std_logic;
	signal And234820_o0 : std_logic;
	signal Or234840_o0 : std_logic;
	signal Nor234860_o0 : std_logic;
	signal And234880_o0 : std_logic;
	signal Or234900_o0 : std_logic;
	signal Or234920_o0 : std_logic;
	signal Or234940_o0 : std_logic;
	signal And234960_o0 : std_logic;
	signal Or234980_o0 : std_logic;
	signal And235000_o0 : std_logic;
	signal Or235020_o0 : std_logic;
	signal And235040_o0 : std_logic;
	signal And235060_o0 : std_logic;
	signal And235080_o0 : std_logic;
	signal Or235100_o0 : std_logic;
	signal Nand235120_o0 : std_logic;
	signal Or235140_o0 : std_logic;
	signal And235160_o0 : std_logic;
	signal And235180_o0 : std_logic;
	signal And235200_o0 : std_logic;
	signal Or235220_o0 : std_logic;
	signal And235240_o0 : std_logic;
	signal And235260_o0 : std_logic;
	signal Or235280_o0 : std_logic;
	signal And235300_o0 : std_logic;
	signal And235320_o0 : std_logic;
	signal Or235340_o0 : std_logic;
	signal And235360_o0 : std_logic;
	signal And235380_o0 : std_logic;
	signal And235400_o0 : std_logic;
	signal And235420_o0 : std_logic;
	signal Or235440_o0 : std_logic;
	signal And235460_o0 : std_logic;
	signal And235480_o0 : std_logic;
	signal And235500_o0 : std_logic;
	signal And235520_o0 : std_logic;
	signal Or235540_o0 : std_logic;
	signal And235560_o0 : std_logic;
	signal And235580_o0 : std_logic;
	signal And235600_o0 : std_logic;
	signal Or235620_o0 : std_logic;
	signal And235640_o0 : std_logic;
	signal And235660_o0 : std_logic;
	signal And235680_o0 : std_logic;
	signal Or235700_o0 : std_logic;
	signal And235720_o0 : std_logic;
	signal And235740_o0 : std_logic;
	signal And235760_o0 : std_logic;
	signal Or235780_o0 : std_logic;
	signal And235800_o0 : std_logic;
	signal Nor235820_o0 : std_logic;
	signal And235840_o0 : std_logic;
	signal Or235860_o0 : std_logic;
	signal And235880_o0 : std_logic;
	signal And235900_o0 : std_logic;
	signal And235920_o0 : std_logic;
	signal Or235940_o0 : std_logic;
	signal And235960_o0 : std_logic;
	signal Or235980_o0 : std_logic;
	signal And236000_o0 : std_logic;
	signal And236020_o0 : std_logic;
	signal And236040_o0 : std_logic;
	signal And236060_o0 : std_logic;
	signal Or236080_o0 : std_logic;
	signal And236100_o0 : std_logic;
	signal And236120_o0 : std_logic;
	signal And236140_o0 : std_logic;
	signal Or236160_o0 : std_logic;
	signal And236180_o0 : std_logic;
	signal And236200_o0 : std_logic;
	signal Or236220_o0 : std_logic;
	signal And236240_o0 : std_logic;
	signal And236260_o0 : std_logic;
	signal Or236280_o0 : std_logic;
	signal And236300_o0 : std_logic;
	signal And236320_o0 : std_logic;
	signal Or236340_o0 : std_logic;
	signal And236360_o0 : std_logic;
	signal Nor236380_o0 : std_logic;
	signal Nor236400_o0 : std_logic;
	signal And236420_o0 : std_logic;
	signal Or236440_o0 : std_logic;
	signal And236460_o0 : std_logic;
	signal Or236480_o0 : std_logic;
	signal And236500_o0 : std_logic;
	signal And236520_o0 : std_logic;
	signal Xor236540_o0 : std_logic;
	signal Or236560_o0 : std_logic;
	signal And236580_o0 : std_logic;
	signal And236600_o0 : std_logic;
	signal Or236620_o0 : std_logic;
	signal And236640_o0 : std_logic;
	signal And236660_o0 : std_logic;
	signal And236680_o0 : std_logic;
	signal And236700_o0 : std_logic;
	signal And236720_o0 : std_logic;
	signal Or236740_o0 : std_logic;
	signal Or236760_o0 : std_logic;
	signal Or236780_o0 : std_logic;
	signal And236800_o0 : std_logic;
	signal And236820_o0 : std_logic;
	signal Nor236840_o0 : std_logic;
	signal And236860_o0 : std_logic;
	signal And236880_o0 : std_logic;
	signal Or236900_o0 : std_logic;
	signal And236920_o0 : std_logic;
	signal And236940_o0 : std_logic;
	signal Or236960_o0 : std_logic;
	signal And236980_o0 : std_logic;
	signal And237000_o0 : std_logic;
	signal Or237020_o0 : std_logic;
	signal And237040_o0 : std_logic;
	signal And237060_o0 : std_logic;
	signal And237080_o0 : std_logic;
	signal And237100_o0 : std_logic;
	signal Or237120_o0 : std_logic;
	signal And237140_o0 : std_logic;
	signal Or237160_o0 : std_logic;
	signal And237180_o0 : std_logic;
	signal And237200_o0 : std_logic;
	signal And237220_o0 : std_logic;
	signal Or237240_o0 : std_logic;
	signal And237260_o0 : std_logic;
	signal And237280_o0 : std_logic;
	signal And237300_o0 : std_logic;
	signal Or237320_o0 : std_logic;
	signal And237340_o0 : std_logic;
	signal And237360_o0 : std_logic;
	signal Or237380_o0 : std_logic;
	signal And237400_o0 : std_logic;
	signal Or237420_o0 : std_logic;
	signal And237440_o0 : std_logic;
	signal And237460_o0 : std_logic;
	signal And237480_o0 : std_logic;
	signal Or237500_o0 : std_logic;
	signal And237520_o0 : std_logic;
	signal And237540_o0 : std_logic;
	signal And237560_o0 : std_logic;
	signal Nor237580_o0 : std_logic;
	signal And237600_o0 : std_logic;
	signal And237620_o0 : std_logic;
	signal And237640_o0 : std_logic;
	signal Or237660_o0 : std_logic;
	signal And237680_o0 : std_logic;
	signal Xor237700_o0 : std_logic;
	signal And237720_o0 : std_logic;
	signal Or237740_o0 : std_logic;
	signal And237760_o0 : std_logic;
	signal Or237780_o0 : std_logic;
	signal And237800_o0 : std_logic;
	signal Or237820_o0 : std_logic;
	signal And237840_o0 : std_logic;
	signal And237860_o0 : std_logic;
	signal And237880_o0 : std_logic;
	signal Or237900_o0 : std_logic;
	signal And237920_o0 : std_logic;
	signal And237940_o0 : std_logic;
	signal And237960_o0 : std_logic;
	signal And237980_o0 : std_logic;
	signal And238000_o0 : std_logic;
	signal Or238020_o0 : std_logic;
	signal And238040_o0 : std_logic;
	signal And238060_o0 : std_logic;
	signal Or238080_o0 : std_logic;
	signal And238100_o0 : std_logic;
	signal Nor238120_o0 : std_logic;
	signal And238140_o0 : std_logic;
	signal And238160_o0 : std_logic;
	signal Or238180_o0 : std_logic;
	signal And238200_o0 : std_logic;
	signal And238220_o0 : std_logic;
	signal And238240_o0 : std_logic;
	signal Or238260_o0 : std_logic;
	signal And238280_o0 : std_logic;
	signal And238300_o0 : std_logic;
	signal Or238320_o0 : std_logic;
	signal And238340_o0 : std_logic;
	signal And238360_o0 : std_logic;
	signal And238380_o0 : std_logic;
	signal Nor238400_o0 : std_logic;
	signal Or238420_o0 : std_logic;
	signal And238440_o0 : std_logic;
	signal And238460_o0 : std_logic;
	signal And238480_o0 : std_logic;
	signal And238500_o0 : std_logic;
	signal Or238520_o0 : std_logic;
	signal And238540_o0 : std_logic;
	signal And238560_o0 : std_logic;
	signal Or238580_o0 : std_logic;
	signal And238600_o0 : std_logic;
	signal And238620_o0 : std_logic;
	signal And238640_o0 : std_logic;
	signal And238660_o0 : std_logic;
	signal Or238680_o0 : std_logic;
	signal And238700_o0 : std_logic;
	signal And238720_o0 : std_logic;
	signal And238740_o0 : std_logic;
	signal Or238760_o0 : std_logic;
	signal And238780_o0 : std_logic;
	signal Or238800_o0 : std_logic;
	signal And238820_o0 : std_logic;
	signal And238840_o0 : std_logic;
	signal And238860_o0 : std_logic;
	signal Or238880_o0 : std_logic;
	signal And238900_o0 : std_logic;
	signal Or238920_o0 : std_logic;
	signal And238940_o0 : std_logic;
	signal Or238960_o0 : std_logic;
	signal And238980_o0 : std_logic;
	signal And239000_o0 : std_logic;
	signal And239020_o0 : std_logic;
	signal Or239040_o0 : std_logic;
	signal Or239060_o0 : std_logic;
	signal Or239080_o0 : std_logic;
	signal And239100_o0 : std_logic;
	signal And239120_o0 : std_logic;
	signal And239140_o0 : std_logic;
	signal Or239160_o0 : std_logic;
	signal Or239180_o0 : std_logic;
	signal And239200_o0 : std_logic;
	signal Xor239220_o0 : std_logic;
	signal And239240_o0 : std_logic;
	signal And239260_o0 : std_logic;
	signal Or239280_o0 : std_logic;
	signal And239300_o0 : std_logic;
	signal And239320_o0 : std_logic;
	signal And239340_o0 : std_logic;
	signal And239360_o0 : std_logic;
	signal Or239380_o0 : std_logic;
	signal And239400_o0 : std_logic;
	signal And239420_o0 : std_logic;
	signal Or239440_o0 : std_logic;
	signal And239460_o0 : std_logic;
	signal Or239480_o0 : std_logic;
	signal And239500_o0 : std_logic;
	signal And239520_o0 : std_logic;
	signal Or239540_o0 : std_logic;
	signal And239560_o0 : std_logic;
	signal And239580_o0 : std_logic;
	signal And239600_o0 : std_logic;
	signal And239620_o0 : std_logic;
	signal And239640_o0 : std_logic;
	signal Or239660_o0 : std_logic;
	signal And239680_o0 : std_logic;
	signal And239700_o0 : std_logic;
	signal Or239720_o0 : std_logic;
	signal And239740_o0 : std_logic;
	signal And239760_o0 : std_logic;
	signal And239780_o0 : std_logic;
	signal Or239800_o0 : std_logic;
	signal And239820_o0 : std_logic;
	signal And239840_o0 : std_logic;
	signal And239860_o0 : std_logic;
	signal And239880_o0 : std_logic;
	signal Or239900_o0 : std_logic;
	signal Or239920_o0 : std_logic;
	signal Or239940_o0 : std_logic;
	signal Or239960_o0 : std_logic;
	signal Or239980_o0 : std_logic;
	signal And240000_o0 : std_logic;
	signal Or240020_o0 : std_logic;
	signal And240040_o0 : std_logic;
	signal And240060_o0 : std_logic;
	signal Or240080_o0 : std_logic;
	signal Or240100_o0 : std_logic;
	signal And240120_o0 : std_logic;
	signal And240140_o0 : std_logic;
	signal And240160_o0 : std_logic;
	signal And240180_o0 : std_logic;
	signal Or240200_o0 : std_logic;
	signal Or240220_o0 : std_logic;
	signal Or240240_o0 : std_logic;
	signal And240260_o0 : std_logic;
	signal And240280_o0 : std_logic;
	signal Or240300_o0 : std_logic;
	signal And240320_o0 : std_logic;
	signal And240340_o0 : std_logic;
	signal And240360_o0 : std_logic;
	signal And240380_o0 : std_logic;
	signal And240400_o0 : std_logic;
	signal And240420_o0 : std_logic;
	signal Or240440_o0 : std_logic;
	signal And240460_o0 : std_logic;
	signal And240480_o0 : std_logic;
	signal Or240500_o0 : std_logic;
	signal And240520_o0 : std_logic;
	signal And240540_o0 : std_logic;
	signal And240560_o0 : std_logic;
	signal And240580_o0 : std_logic;
	signal Or240600_o0 : std_logic;
	signal And240620_o0 : std_logic;
	signal And240640_o0 : std_logic;
	signal And240660_o0 : std_logic;
	signal Or240680_o0 : std_logic;
	signal Or240700_o0 : std_logic;
	signal And240720_o0 : std_logic;
	signal And240740_o0 : std_logic;
	signal Nor240760_o0 : std_logic;
	signal And240780_o0 : std_logic;
	signal Or240800_o0 : std_logic;
	signal And240820_o0 : std_logic;
	signal And240840_o0 : std_logic;
	signal Or240860_o0 : std_logic;
	signal And240880_o0 : std_logic;
	signal And240900_o0 : std_logic;
	signal And240920_o0 : std_logic;
	signal Or240940_o0 : std_logic;
	signal And240960_o0 : std_logic;
	signal Or240980_o0 : std_logic;
	signal And241000_o0 : std_logic;
	signal Or241020_o0 : std_logic;
	signal And241040_o0 : std_logic;
	signal And241060_o0 : std_logic;
	signal And241080_o0 : std_logic;
	signal Or241100_o0 : std_logic;
	signal And241120_o0 : std_logic;
	signal Or241140_o0 : std_logic;
	signal And241160_o0 : std_logic;
	signal And241180_o0 : std_logic;
	signal Or241200_o0 : std_logic;
	signal And241220_o0 : std_logic;
	signal And241240_o0 : std_logic;
	signal Or241260_o0 : std_logic;
	signal And241280_o0 : std_logic;
	signal And241300_o0 : std_logic;
	signal And241320_o0 : std_logic;
	signal Or241340_o0 : std_logic;
	signal And241360_o0 : std_logic;
	signal And241380_o0 : std_logic;
	signal Or241400_o0 : std_logic;
	signal And241420_o0 : std_logic;
	signal And241440_o0 : std_logic;
	signal And241460_o0 : std_logic;
	signal And241480_o0 : std_logic;
	signal And241500_o0 : std_logic;
	signal Or241520_o0 : std_logic;
	signal And241540_o0 : std_logic;
	signal And241560_o0 : std_logic;
	signal And241580_o0 : std_logic;
	signal And241600_o0 : std_logic;
	signal And241620_o0 : std_logic;
	signal Or241640_o0 : std_logic;
	signal And241660_o0 : std_logic;
	signal Or241680_o0 : std_logic;
	signal And241700_o0 : std_logic;
	signal And241720_o0 : std_logic;
	signal Or241740_o0 : std_logic;
	signal And241760_o0 : std_logic;
	signal Or241780_o0 : std_logic;
	signal And241800_o0 : std_logic;
	signal Or241820_o0 : std_logic;
	signal And241840_o0 : std_logic;
	signal Or241860_o0 : std_logic;
	signal And241880_o0 : std_logic;
	signal And241900_o0 : std_logic;
	signal Or241920_o0 : std_logic;
	signal And241940_o0 : std_logic;
	signal Or241960_o0 : std_logic;
	signal And241980_o0 : std_logic;
	signal And242000_o0 : std_logic;
	signal And242020_o0 : std_logic;
	signal And242040_o0 : std_logic;
	signal Or242060_o0 : std_logic;
	signal And242080_o0 : std_logic;
	signal And242100_o0 : std_logic;
	signal And242120_o0 : std_logic;
	signal Or242140_o0 : std_logic;
	signal And242160_o0 : std_logic;
	signal And242180_o0 : std_logic;
	signal And242200_o0 : std_logic;
	signal Or242220_o0 : std_logic;
	signal And242240_o0 : std_logic;
	signal And242260_o0 : std_logic;
	signal And242280_o0 : std_logic;
	signal And242300_o0 : std_logic;
	signal Or242320_o0 : std_logic;
	signal And242340_o0 : std_logic;
	signal And242360_o0 : std_logic;
	signal And242380_o0 : std_logic;
	signal And242400_o0 : std_logic;
	signal Or242420_o0 : std_logic;
	signal And242440_o0 : std_logic;
	signal And242460_o0 : std_logic;
	signal And242480_o0 : std_logic;
	signal And242500_o0 : std_logic;
	signal Or242520_o0 : std_logic;
	signal And242540_o0 : std_logic;
	signal And242560_o0 : std_logic;
	signal And242580_o0 : std_logic;
	signal Or242600_o0 : std_logic;
	signal And242620_o0 : std_logic;
	signal And242640_o0 : std_logic;
	signal Or242660_o0 : std_logic;
	signal And242680_o0 : std_logic;
	signal Or242700_o0 : std_logic;
	signal And242720_o0 : std_logic;
	signal And242740_o0 : std_logic;
	signal Or242760_o0 : std_logic;
	signal And242780_o0 : std_logic;
	signal And242800_o0 : std_logic;
	signal And242820_o0 : std_logic;
	signal Or242840_o0 : std_logic;
	signal And242860_o0 : std_logic;
	signal And242880_o0 : std_logic;
	signal Or242900_o0 : std_logic;
	signal And242920_o0 : std_logic;
	signal And242940_o0 : std_logic;
	signal And242960_o0 : std_logic;
	signal Or242980_o0 : std_logic;
	signal And243000_o0 : std_logic;
	signal And243020_o0 : std_logic;
	signal And243040_o0 : std_logic;
	signal And243060_o0 : std_logic;
	signal Or243080_o0 : std_logic;
	signal And243100_o0 : std_logic;
	signal And243120_o0 : std_logic;
	signal Or243140_o0 : std_logic;
	signal And243160_o0 : std_logic;
	signal Or243180_o0 : std_logic;
	signal And243200_o0 : std_logic;
	signal And243220_o0 : std_logic;
	signal Or243240_o0 : std_logic;
	signal And243260_o0 : std_logic;
	signal Or243280_o0 : std_logic;
	signal And243300_o0 : std_logic;
	signal And243320_o0 : std_logic;
	signal And243340_o0 : std_logic;
	signal And243360_o0 : std_logic;
	signal Or243380_o0 : std_logic;
	signal And243400_o0 : std_logic;
	signal Nor243420_o0 : std_logic;
	signal Or243440_o0 : std_logic;
	signal And243460_o0 : std_logic;
	signal And243480_o0 : std_logic;
	signal Or243500_o0 : std_logic;
	signal And243520_o0 : std_logic;
	signal And243540_o0 : std_logic;
	signal And243560_o0 : std_logic;
	signal Or243580_o0 : std_logic;
	signal And243600_o0 : std_logic;
	signal And243620_o0 : std_logic;
	signal Or243640_o0 : std_logic;
	signal And243660_o0 : std_logic;
	signal And243680_o0 : std_logic;
	signal Or243700_o0 : std_logic;
	signal And243720_o0 : std_logic;
	signal Or243740_o0 : std_logic;
	signal Or243760_o0 : std_logic;
	signal And243780_o0 : std_logic;
	signal Or243800_o0 : std_logic;
	signal And243820_o0 : std_logic;
	signal And243840_o0 : std_logic;
	signal And243860_o0 : std_logic;
	signal And243880_o0 : std_logic;
	signal Or243900_o0 : std_logic;
	signal Or243920_o0 : std_logic;
	signal And243940_o0 : std_logic;
	signal And243960_o0 : std_logic;
	signal And243980_o0 : std_logic;
	signal And244000_o0 : std_logic;
	signal Or244020_o0 : std_logic;
	signal And244040_o0 : std_logic;
	signal Or244060_o0 : std_logic;
	signal And244080_o0 : std_logic;
	signal Or244100_o0 : std_logic;
	signal And244120_o0 : std_logic;
	signal And244140_o0 : std_logic;
	signal Or244160_o0 : std_logic;
	signal And244180_o0 : std_logic;
	signal Or244200_o0 : std_logic;
	signal And244220_o0 : std_logic;
	signal Or244240_o0 : std_logic;
	signal Or244260_o0 : std_logic;
	signal And244280_o0 : std_logic;
	signal Or244300_o0 : std_logic;
	signal And244320_o0 : std_logic;
	signal And244340_o0 : std_logic;
	signal And244360_o0 : std_logic;
	signal Or244380_o0 : std_logic;
	signal And244400_o0 : std_logic;
	signal And244420_o0 : std_logic;
	signal Or244440_o0 : std_logic;
	signal And244460_o0 : std_logic;
	signal And244480_o0 : std_logic;
	signal Or244500_o0 : std_logic;
	signal Or244520_o0 : std_logic;
	signal Or244540_o0 : std_logic;
	signal Or244560_o0 : std_logic;
	signal And244580_o0 : std_logic;
	signal And244600_o0 : std_logic;
	signal Or244620_o0 : std_logic;
	signal And244640_o0 : std_logic;
	signal And244660_o0 : std_logic;
	signal Or244680_o0 : std_logic;
	signal And244700_o0 : std_logic;
	signal Or244720_o0 : std_logic;
	signal And244740_o0 : std_logic;
	signal Or244760_o0 : std_logic;
	signal And244780_o0 : std_logic;
	signal And244800_o0 : std_logic;
	signal And244820_o0 : std_logic;
	signal And244840_o0 : std_logic;
	signal And244860_o0 : std_logic;
	signal Or244880_o0 : std_logic;
	signal And244900_o0 : std_logic;
	signal Or244920_o0 : std_logic;
	signal Or244940_o0 : std_logic;
	signal Or244960_o0 : std_logic;
	signal Or244980_o0 : std_logic;
	signal And245000_o0 : std_logic;
	signal Or245020_o0 : std_logic;
	signal And245040_o0 : std_logic;
	signal Or245060_o0 : std_logic;
	signal And245080_o0 : std_logic;
	signal And245100_o0 : std_logic;
	signal And245120_o0 : std_logic;
	signal And245140_o0 : std_logic;
	signal Or245160_o0 : std_logic;
	signal And245180_o0 : std_logic;
	signal And245200_o0 : std_logic;
	signal And245220_o0 : std_logic;
	signal And245240_o0 : std_logic;
	signal And245260_o0 : std_logic;
	signal And245280_o0 : std_logic;
	signal And245300_o0 : std_logic;
	signal Or245320_o0 : std_logic;
	signal And245340_o0 : std_logic;
	signal Or245360_o0 : std_logic;
	signal And245380_o0 : std_logic;
	signal Or245400_o0 : std_logic;
	signal Or245420_o0 : std_logic;
	signal Or245440_o0 : std_logic;
	signal And245460_o0 : std_logic;
	signal Or245480_o0 : std_logic;
	signal And245500_o0 : std_logic;
	signal Or245520_o0 : std_logic;
	signal And245540_o0 : std_logic;
	signal Nand245560_o0 : std_logic;
	signal Or245580_o0 : std_logic;
	signal And245600_o0 : std_logic;
	signal And245620_o0 : std_logic;
	signal Or245640_o0 : std_logic;
	signal And245660_o0 : std_logic;
	signal Xor245680_o0 : std_logic;
	signal And245700_o0 : std_logic;
	signal And245720_o0 : std_logic;
	signal And245740_o0 : std_logic;
	signal Or245760_o0 : std_logic;
	signal Or245780_o0 : std_logic;
	signal Or245800_o0 : std_logic;
	signal And245820_o0 : std_logic;
	signal And245840_o0 : std_logic;
	signal Or245860_o0 : std_logic;
	signal And245880_o0 : std_logic;
	signal Or245900_o0 : std_logic;
	signal Or245920_o0 : std_logic;
	signal And245940_o0 : std_logic;
	signal Or245960_o0 : std_logic;
	signal And245980_o0 : std_logic;
	signal Xor246000_o0 : std_logic;
	signal Not46020_o0 : std_logic;
	signal Or246040_o0 : std_logic;
	signal And246060_o0 : std_logic;
	signal Or246080_o0 : std_logic;
	signal Or246100_o0 : std_logic;
	signal And246120_o0 : std_logic;
	signal Or246140_o0 : std_logic;
	signal And246160_o0 : std_logic;
	signal And246180_o0 : std_logic;
	signal And246200_o0 : std_logic;
	signal Or246220_o0 : std_logic;
	signal And246240_o0 : std_logic;
	signal And246260_o0 : std_logic;
	signal And246280_o0 : std_logic;
	signal Or246300_o0 : std_logic;
	signal And246320_o0 : std_logic;
	signal And246340_o0 : std_logic;
	signal Or246360_o0 : std_logic;
	signal And246380_o0 : std_logic;
	signal And246400_o0 : std_logic;
	signal Or246420_o0 : std_logic;
	signal And246440_o0 : std_logic;
	signal Or246460_o0 : std_logic;
	signal And246480_o0 : std_logic;
	signal Or246500_o0 : std_logic;
	signal And246520_o0 : std_logic;
	signal And246540_o0 : std_logic;
	signal Or246560_o0 : std_logic;
	signal And246580_o0 : std_logic;
	signal Or246600_o0 : std_logic;
	signal And246620_o0 : std_logic;
	signal And246640_o0 : std_logic;
	signal And246660_o0 : std_logic;
	signal And246680_o0 : std_logic;
	signal Or246700_o0 : std_logic;
	signal And246720_o0 : std_logic;
	signal Or246740_o0 : std_logic;
	signal And246760_o0 : std_logic;
	signal And246780_o0 : std_logic;
	signal And246800_o0 : std_logic;
	signal Or246820_o0 : std_logic;
	signal And246840_o0 : std_logic;
	signal And246860_o0 : std_logic;
	signal Or246880_o0 : std_logic;
	signal And246900_o0 : std_logic;
	signal And246920_o0 : std_logic;
	signal And246940_o0 : std_logic;
	signal And246960_o0 : std_logic;
	signal And246980_o0 : std_logic;
	signal Or247000_o0 : std_logic;
	signal And247020_o0 : std_logic;
	signal And247040_o0 : std_logic;
	signal And247060_o0 : std_logic;
	signal And247080_o0 : std_logic;
	signal Or247100_o0 : std_logic;
	signal Or247120_o0 : std_logic;
	signal Or247140_o0 : std_logic;
	signal Or247160_o0 : std_logic;
	signal And247180_o0 : std_logic;
	signal Or247200_o0 : std_logic;
	signal And247220_o0 : std_logic;
	signal And247240_o0 : std_logic;
	signal Or247260_o0 : std_logic;
	signal And247280_o0 : std_logic;
	signal And247300_o0 : std_logic;
	signal Or247320_o0 : std_logic;
	signal And247340_o0 : std_logic;
	signal Or247360_o0 : std_logic;
	signal And247380_o0 : std_logic;
	signal And247400_o0 : std_logic;
	signal And247420_o0 : std_logic;
	signal Or247440_o0 : std_logic;
	signal And247460_o0 : std_logic;
	signal Or247480_o0 : std_logic;
	signal And247500_o0 : std_logic;
	signal Or247520_o0 : std_logic;
	signal And247540_o0 : std_logic;
	signal And247560_o0 : std_logic;
	signal And247580_o0 : std_logic;
	signal And247600_o0 : std_logic;
	signal Or247620_o0 : std_logic;
	signal And247640_o0 : std_logic;
	signal And247660_o0 : std_logic;
	signal Nor247680_o0 : std_logic;
	signal Or247700_o0 : std_logic;
	signal And247720_o0 : std_logic;
	signal And247740_o0 : std_logic;
	signal Or247760_o0 : std_logic;
	signal And247780_o0 : std_logic;
	signal And247800_o0 : std_logic;
	signal And247820_o0 : std_logic;
	signal Or247840_o0 : std_logic;
	signal And247860_o0 : std_logic;
	signal Not47880_o0 : std_logic;
	signal Nor247900_o0 : std_logic;
	signal Or247920_o0 : std_logic;
	signal And247940_o0 : std_logic;
	signal Or247960_o0 : std_logic;
	signal And247980_o0 : std_logic;
	signal And248000_o0 : std_logic;
	signal And248020_o0 : std_logic;
	signal And248040_o0 : std_logic;
	signal Or248060_o0 : std_logic;
	signal And248080_o0 : std_logic;
	signal Or248100_o0 : std_logic;
	signal Or248120_o0 : std_logic;
	signal And248140_o0 : std_logic;
	signal And248160_o0 : std_logic;
	signal And248180_o0 : std_logic;
	signal And248200_o0 : std_logic;
	signal Or248220_o0 : std_logic;
	signal And248240_o0 : std_logic;
	signal And248260_o0 : std_logic;
	signal And248280_o0 : std_logic;
	signal And248300_o0 : std_logic;
	signal And248320_o0 : std_logic;
	signal And248340_o0 : std_logic;
	signal And248360_o0 : std_logic;
	signal Or248380_o0 : std_logic;
	signal And248400_o0 : std_logic;
	signal And248420_o0 : std_logic;
	signal And248440_o0 : std_logic;
	signal And248460_o0 : std_logic;
	signal Or248480_o0 : std_logic;
	signal And248500_o0 : std_logic;
	signal And248520_o0 : std_logic;
	signal And248540_o0 : std_logic;
	signal And248560_o0 : std_logic;
	signal Or248580_o0 : std_logic;
	signal And248600_o0 : std_logic;
	signal Or248620_o0 : std_logic;
	signal And248640_o0 : std_logic;
	signal Nor248660_o0 : std_logic;
	signal And248680_o0 : std_logic;
	signal And248700_o0 : std_logic;
	signal And248720_o0 : std_logic;
	signal Or248740_o0 : std_logic;
	signal And248760_o0 : std_logic;
	signal Or248780_o0 : std_logic;
	signal And248800_o0 : std_logic;
	signal Or248820_o0 : std_logic;
	signal And248840_o0 : std_logic;
	signal And248860_o0 : std_logic;
	signal Or248880_o0 : std_logic;
	signal And248900_o0 : std_logic;
	signal And248920_o0 : std_logic;
	signal And248940_o0 : std_logic;
	signal Or248960_o0 : std_logic;
	signal And248980_o0 : std_logic;
	signal And249000_o0 : std_logic;
	signal And249020_o0 : std_logic;
	signal And249040_o0 : std_logic;
	signal Or249060_o0 : std_logic;
	signal And249080_o0 : std_logic;
	signal Or249100_o0 : std_logic;
	signal And249120_o0 : std_logic;
	signal Or249140_o0 : std_logic;
	signal And249160_o0 : std_logic;
	signal Or249180_o0 : std_logic;
	signal And249200_o0 : std_logic;
	signal Or249220_o0 : std_logic;
	signal And249240_o0 : std_logic;
	signal Or249260_o0 : std_logic;
	signal And249280_o0 : std_logic;
	signal And249300_o0 : std_logic;
	signal Or249320_o0 : std_logic;
	signal And249340_o0 : std_logic;
	signal Or249360_o0 : std_logic;
	signal Or249380_o0 : std_logic;
	signal And249400_o0 : std_logic;
	signal Or249420_o0 : std_logic;
	signal And249440_o0 : std_logic;
	signal And249460_o0 : std_logic;
	signal And249480_o0 : std_logic;
	signal Or249500_o0 : std_logic;
	signal Or249520_o0 : std_logic;
	signal Or249540_o0 : std_logic;
	signal Or249560_o0 : std_logic;
	signal And249580_o0 : std_logic;
	signal Or249600_o0 : std_logic;
	signal And249620_o0 : std_logic;
	signal And249640_o0 : std_logic;
	signal Or249660_o0 : std_logic;
	signal Or249680_o0 : std_logic;
	signal And249700_o0 : std_logic;
	signal Or249720_o0 : std_logic;
	signal And249740_o0 : std_logic;
	signal Or249760_o0 : std_logic;
	signal And249780_o0 : std_logic;
	signal Or249800_o0 : std_logic;
	signal And249820_o0 : std_logic;
	signal Or249840_o0 : std_logic;
	signal And249860_o0 : std_logic;
	signal And249880_o0 : std_logic;
	signal And249900_o0 : std_logic;
	signal Or249920_o0 : std_logic;
	signal And249940_o0 : std_logic;
	signal And249960_o0 : std_logic;
	signal And249980_o0 : std_logic;
	signal Or250000_o0 : std_logic;
	signal Or250020_o0 : std_logic;
	signal Or250040_o0 : std_logic;
	signal And250060_o0 : std_logic;
	signal Or250080_o0 : std_logic;
	signal And250100_o0 : std_logic;
	signal And250120_o0 : std_logic;
	signal Or250140_o0 : std_logic;
	signal And250160_o0 : std_logic;
	signal And250180_o0 : std_logic;
	signal Or250200_o0 : std_logic;
	signal And250220_o0 : std_logic;
	signal Or250240_o0 : std_logic;
	signal And250260_o0 : std_logic;
	signal And250280_o0 : std_logic;
	signal And250300_o0 : std_logic;
	signal Nor250320_o0 : std_logic;
	signal And250340_o0 : std_logic;
	signal And250360_o0 : std_logic;
	signal Or250380_o0 : std_logic;
	signal Or250400_o0 : std_logic;
	signal And250420_o0 : std_logic;
	signal Or250440_o0 : std_logic;
	signal And250460_o0 : std_logic;
	signal And250480_o0 : std_logic;
	signal And250500_o0 : std_logic;
	signal Or250520_o0 : std_logic;
	signal Or250540_o0 : std_logic;
	signal Or250560_o0 : std_logic;
	signal Or250580_o0 : std_logic;
	signal And250600_o0 : std_logic;
	signal Or250620_o0 : std_logic;
	signal Or250640_o0 : std_logic;
	signal And250660_o0 : std_logic;
	signal And250680_o0 : std_logic;
	signal Or250700_o0 : std_logic;
	signal And250720_o0 : std_logic;
	signal And250740_o0 : std_logic;
	signal Or250760_o0 : std_logic;
	signal And250780_o0 : std_logic;
	signal And250800_o0 : std_logic;
	signal Or250820_o0 : std_logic;
	signal And250840_o0 : std_logic;
	signal Or250860_o0 : std_logic;
	signal And250880_o0 : std_logic;
	signal And250900_o0 : std_logic;
	signal Or250920_o0 : std_logic;
	signal Or250940_o0 : std_logic;
	signal Or250960_o0 : std_logic;
	signal Or250980_o0 : std_logic;
	signal And251000_o0 : std_logic;
	signal Or251020_o0 : std_logic;
	signal And251040_o0 : std_logic;
	signal Or251060_o0 : std_logic;
	signal And251080_o0 : std_logic;
	signal And251100_o0 : std_logic;
	signal And251120_o0 : std_logic;
	signal And251140_o0 : std_logic;
	signal And251160_o0 : std_logic;
	signal And251180_o0 : std_logic;
	signal Or251200_o0 : std_logic;
	signal And251220_o0 : std_logic;
	signal Or251240_o0 : std_logic;
	signal And251260_o0 : std_logic;
	signal Or251280_o0 : std_logic;
	signal And251300_o0 : std_logic;
	signal Or251320_o0 : std_logic;
	signal Or251340_o0 : std_logic;
	signal And251360_o0 : std_logic;
	signal Or251380_o0 : std_logic;
	signal And251400_o0 : std_logic;
	signal Or251420_o0 : std_logic;
	signal Or251440_o0 : std_logic;
	signal And251460_o0 : std_logic;
	signal Or251480_o0 : std_logic;
	signal And251500_o0 : std_logic;
	signal Or251520_o0 : std_logic;
	signal And251540_o0 : std_logic;
	signal Or251560_o0 : std_logic;
	signal And251580_o0 : std_logic;
	signal Or251600_o0 : std_logic;
	signal And251620_o0 : std_logic;
	signal Or251640_o0 : std_logic;
	signal And251660_o0 : std_logic;
	signal Or251680_o0 : std_logic;
	signal And251700_o0 : std_logic;
	signal Or251720_o0 : std_logic;
	signal And251740_o0 : std_logic;
	signal Or251760_o0 : std_logic;
	signal And251780_o0 : std_logic;
	signal Or251800_o0 : std_logic;
	signal And251820_o0 : std_logic;
	signal Or251840_o0 : std_logic;
	signal Xor251860_o0 : std_logic;
	signal Or251880_o0 : std_logic;
	signal And251900_o0 : std_logic;
	signal And251920_o0 : std_logic;
	signal And251940_o0 : std_logic;
	signal Or251960_o0 : std_logic;
	signal And251980_o0 : std_logic;
	signal And252000_o0 : std_logic;
	signal Nor252020_o0 : std_logic;
	signal And252040_o0 : std_logic;
	signal And252060_o0 : std_logic;
	signal And252080_o0 : std_logic;
	signal And252100_o0 : std_logic;
	signal Or252120_o0 : std_logic;
	signal And252140_o0 : std_logic;
	signal Or252160_o0 : std_logic;
	signal And252180_o0 : std_logic;
	signal Or252200_o0 : std_logic;
	signal And252220_o0 : std_logic;
	signal Or252240_o0 : std_logic;
	signal And252260_o0 : std_logic;
	signal Or252280_o0 : std_logic;
	signal Or252300_o0 : std_logic;
	signal And252320_o0 : std_logic;
	signal Or252340_o0 : std_logic;
	signal And252360_o0 : std_logic;
	signal Or252380_o0 : std_logic;
	signal Or252400_o0 : std_logic;
	signal And252420_o0 : std_logic;
	signal And252440_o0 : std_logic;
	signal Or252460_o0 : std_logic;
	signal And252480_o0 : std_logic;
	signal And252500_o0 : std_logic;
	signal And252520_o0 : std_logic;
	signal Or252540_o0 : std_logic;
	signal And252560_o0 : std_logic;
	signal And252580_o0 : std_logic;
	signal And252600_o0 : std_logic;
	signal Or252620_o0 : std_logic;
	signal And252640_o0 : std_logic;
	signal And252660_o0 : std_logic;
	signal And252680_o0 : std_logic;
	signal Or252700_o0 : std_logic;
	signal And252720_o0 : std_logic;
	signal And252740_o0 : std_logic;
	signal And252760_o0 : std_logic;
	signal Or252780_o0 : std_logic;
	signal And252800_o0 : std_logic;
	signal And252820_o0 : std_logic;
	signal And252840_o0 : std_logic;
	signal Or252860_o0 : std_logic;
	signal And252880_o0 : std_logic;
	signal And252900_o0 : std_logic;
	signal And252920_o0 : std_logic;
	signal And252940_o0 : std_logic;
	signal Or252960_o0 : std_logic;
	signal And252980_o0 : std_logic;
	signal And253000_o0 : std_logic;
	signal And253020_o0 : std_logic;
	signal Or253040_o0 : std_logic;
	signal And253060_o0 : std_logic;
	signal Or253080_o0 : std_logic;
	signal And253100_o0 : std_logic;
	signal Or253120_o0 : std_logic;
	signal And253140_o0 : std_logic;
	signal Or253160_o0 : std_logic;
	signal And253180_o0 : std_logic;
	signal Or253200_o0 : std_logic;
	signal And253220_o0 : std_logic;
	signal Or253240_o0 : std_logic;
	signal And253260_o0 : std_logic;
	signal And253280_o0 : std_logic;
	signal And253300_o0 : std_logic;
	signal Or253320_o0 : std_logic;
	signal And253340_o0 : std_logic;
	signal Or253360_o0 : std_logic;
	signal And253380_o0 : std_logic;
	signal Or253400_o0 : std_logic;
	signal And253420_o0 : std_logic;
	signal Or253440_o0 : std_logic;
	signal Or253460_o0 : std_logic;
	signal And253480_o0 : std_logic;
	signal Or253500_o0 : std_logic;
	signal And253520_o0 : std_logic;
	signal Or253540_o0 : std_logic;
	signal And253560_o0 : std_logic;
	signal Or253580_o0 : std_logic;
	signal And253600_o0 : std_logic;
	signal Or253620_o0 : std_logic;
	signal And253640_o0 : std_logic;
	signal Or253660_o0 : std_logic;
	signal And253680_o0 : std_logic;
	signal Or253700_o0 : std_logic;
	signal And253720_o0 : std_logic;
	signal Or253740_o0 : std_logic;
	signal And253760_o0 : std_logic;
	signal Or253780_o0 : std_logic;
	signal And253800_o0 : std_logic;
	signal Or253820_o0 : std_logic;
	signal And253840_o0 : std_logic;
	signal And253860_o0 : std_logic;
	signal Or253880_o0 : std_logic;
	signal And253900_o0 : std_logic;
	signal Or253920_o0 : std_logic;
	signal And253940_o0 : std_logic;
	signal And253960_o0 : std_logic;
	signal And253980_o0 : std_logic;
	signal And254000_o0 : std_logic;
	signal And254020_o0 : std_logic;
	signal And254040_o0 : std_logic;
	signal And254060_o0 : std_logic;
	signal Or254080_o0 : std_logic;
	signal And254100_o0 : std_logic;
	signal Or254120_o0 : std_logic;
	signal And254140_o0 : std_logic;
	signal And254160_o0 : std_logic;
	signal Or254180_o0 : std_logic;
	signal And254200_o0 : std_logic;
	signal And254220_o0 : std_logic;
	signal And254240_o0 : std_logic;
	signal And254260_o0 : std_logic;
	signal Or254280_o0 : std_logic;
	signal And254300_o0 : std_logic;
	signal And254320_o0 : std_logic;
	signal And254340_o0 : std_logic;
	signal Or254360_o0 : std_logic;
	signal And254380_o0 : std_logic;
	signal And254400_o0 : std_logic;
	signal And254420_o0 : std_logic;
	signal Or254440_o0 : std_logic;
	signal And254460_o0 : std_logic;
	signal And254480_o0 : std_logic;
	signal And254500_o0 : std_logic;
	signal Or254520_o0 : std_logic;
	signal And254540_o0 : std_logic;
	signal And254560_o0 : std_logic;
	signal And254580_o0 : std_logic;
	signal And254600_o0 : std_logic;
	signal And254620_o0 : std_logic;
	signal And254640_o0 : std_logic;
	signal And254660_o0 : std_logic;
	signal Or254680_o0 : std_logic;
	signal And254700_o0 : std_logic;
	signal And254720_o0 : std_logic;
	signal And254740_o0 : std_logic;
	signal And254760_o0 : std_logic;
	signal Or254780_o0 : std_logic;
	signal And254800_o0 : std_logic;
	signal And254820_o0 : std_logic;
	signal Nor254840_o0 : std_logic;
	signal And254860_o0 : std_logic;
	signal Or254880_o0 : std_logic;
	signal And254900_o0 : std_logic;
	signal Or254920_o0 : std_logic;
	signal And254940_o0 : std_logic;
	signal Or254960_o0 : std_logic;
	signal And254980_o0 : std_logic;
	signal And255000_o0 : std_logic;
	signal And255020_o0 : std_logic;
	signal And255040_o0 : std_logic;
	signal And255060_o0 : std_logic;
	signal Or255080_o0 : std_logic;
	signal And255100_o0 : std_logic;
	signal And255120_o0 : std_logic;
	signal And255140_o0 : std_logic;
	signal And255160_o0 : std_logic;
	signal And255180_o0 : std_logic;
	signal Or255200_o0 : std_logic;
	signal And255220_o0 : std_logic;
	signal And255240_o0 : std_logic;
	signal And255260_o0 : std_logic;
	signal Or255280_o0 : std_logic;
	signal And255300_o0 : std_logic;
	signal And255320_o0 : std_logic;
	signal And255340_o0 : std_logic;
	signal And255360_o0 : std_logic;
	signal And255380_o0 : std_logic;
	signal Or255400_o0 : std_logic;
	signal And255420_o0 : std_logic;
	signal And255440_o0 : std_logic;
	signal And255460_o0 : std_logic;
	signal And255480_o0 : std_logic;
	signal And255500_o0 : std_logic;
	signal Or255520_o0 : std_logic;
	signal Nor255540_o0 : std_logic;
	signal And255560_o0 : std_logic;
	signal And255580_o0 : std_logic;
	signal And255600_o0 : std_logic;
	signal And255620_o0 : std_logic;
	signal And255640_o0 : std_logic;
	signal And255660_o0 : std_logic;
	signal And255680_o0 : std_logic;
	signal Or255700_o0 : std_logic;
	signal And255720_o0 : std_logic;
	signal And255740_o0 : std_logic;
	signal And255760_o0 : std_logic;
	signal Or255780_o0 : std_logic;
	signal And255800_o0 : std_logic;
	signal And255820_o0 : std_logic;
	signal And255840_o0 : std_logic;
	signal Or255860_o0 : std_logic;
	signal And255880_o0 : std_logic;
	signal And255900_o0 : std_logic;
	signal And255920_o0 : std_logic;
	signal Or255940_o0 : std_logic;
	signal And255960_o0 : std_logic;
	signal And255980_o0 : std_logic;
	signal And256000_o0 : std_logic;
	signal Or256020_o0 : std_logic;
	signal And256040_o0 : std_logic;
	signal And256060_o0 : std_logic;
	signal And256080_o0 : std_logic;
	signal And256100_o0 : std_logic;
	signal Or256120_o0 : std_logic;
	signal And256140_o0 : std_logic;
	signal And256160_o0 : std_logic;
	signal And256180_o0 : std_logic;
	signal And256200_o0 : std_logic;
	signal Or256220_o0 : std_logic;
	signal And256240_o0 : std_logic;
	signal And256260_o0 : std_logic;
	signal And256280_o0 : std_logic;
	signal And256300_o0 : std_logic;
	signal And256320_o0 : std_logic;
	signal And256340_o0 : std_logic;
	signal Or256360_o0 : std_logic;
	signal And256380_o0 : std_logic;
	signal And256400_o0 : std_logic;
	signal And256420_o0 : std_logic;
	signal Or256440_o0 : std_logic;
	signal And256460_o0 : std_logic;
	signal And256480_o0 : std_logic;
	signal And256500_o0 : std_logic;
	signal And256520_o0 : std_logic;
	signal Or256540_o0 : std_logic;
	signal And256560_o0 : std_logic;
	signal And256580_o0 : std_logic;
	signal And256600_o0 : std_logic;
	signal And256620_o0 : std_logic;
	signal Or256640_o0 : std_logic;
	signal And256660_o0 : std_logic;
	signal And256680_o0 : std_logic;
	signal And256700_o0 : std_logic;
	signal And256720_o0 : std_logic;
	signal And256740_o0 : std_logic;
	signal Or256760_o0 : std_logic;
	signal And256780_o0 : std_logic;
	signal And256800_o0 : std_logic;
	signal And256820_o0 : std_logic;
	signal And256840_o0 : std_logic;
	signal And256860_o0 : std_logic;
	signal Nor256880_o0 : std_logic;
	signal And256900_o0 : std_logic;
	signal Or256920_o0 : std_logic;
	signal And256940_o0 : std_logic;
	signal And256960_o0 : std_logic;
	signal And256980_o0 : std_logic;
	signal Or257000_o0 : std_logic;
	signal And257020_o0 : std_logic;
	signal And257040_o0 : std_logic;
	signal Or257060_o0 : std_logic;
	signal And257080_o0 : std_logic;
	signal And257100_o0 : std_logic;
	signal Or257120_o0 : std_logic;
	signal And257140_o0 : std_logic;
	signal And257160_o0 : std_logic;
	signal And257180_o0 : std_logic;
	signal Or257200_o0 : std_logic;
	signal And257220_o0 : std_logic;
	signal Nor257240_o0 : std_logic;
	signal And257260_o0 : std_logic;
	signal Or257280_o0 : std_logic;
	signal And257300_o0 : std_logic;
	signal And257320_o0 : std_logic;
	signal And257340_o0 : std_logic;
	signal And257360_o0 : std_logic;
	signal Or257380_o0 : std_logic;
	signal And257400_o0 : std_logic;
	signal And257420_o0 : std_logic;
	signal And257440_o0 : std_logic;
	signal And257460_o0 : std_logic;
	signal And257480_o0 : std_logic;
	signal Or257500_o0 : std_logic;
	signal And257520_o0 : std_logic;
	signal Or257540_o0 : std_logic;
	signal And257560_o0 : std_logic;
	signal And257580_o0 : std_logic;
	signal And257600_o0 : std_logic;
	signal And257620_o0 : std_logic;
	signal Or257640_o0 : std_logic;
	signal Or257660_o0 : std_logic;
	signal And257680_o0 : std_logic;
	signal And257700_o0 : std_logic;
	signal And257720_o0 : std_logic;
	signal Or257740_o0 : std_logic;
	signal And257760_o0 : std_logic;
	signal Or257780_o0 : std_logic;
	signal And257800_o0 : std_logic;
	signal Or257820_o0 : std_logic;
	signal And257840_o0 : std_logic;
	signal And257860_o0 : std_logic;
	signal And257880_o0 : std_logic;
	signal Or257900_o0 : std_logic;
	signal And257920_o0 : std_logic;
	signal And257940_o0 : std_logic;
	signal And257960_o0 : std_logic;
	signal And257980_o0 : std_logic;
	signal Or258000_o0 : std_logic;
	signal And258020_o0 : std_logic;
	signal Or258040_o0 : std_logic;
	signal And258060_o0 : std_logic;
	signal And258080_o0 : std_logic;
	signal And258100_o0 : std_logic;
	signal Or258120_o0 : std_logic;
	signal And258140_o0 : std_logic;
	signal And258160_o0 : std_logic;
	signal And258180_o0 : std_logic;
	signal And258200_o0 : std_logic;
	signal Or258220_o0 : std_logic;
	signal And258240_o0 : std_logic;
	signal And258260_o0 : std_logic;
	signal Or258280_o0 : std_logic;
	signal And258300_o0 : std_logic;
	signal Or258320_o0 : std_logic;
	signal And258340_o0 : std_logic;
	signal And258360_o0 : std_logic;
	signal Nor258380_o0 : std_logic;
	signal And258400_o0 : std_logic;
	signal Or258420_o0 : std_logic;
	signal And258440_o0 : std_logic;
	signal And258460_o0 : std_logic;
	signal And258480_o0 : std_logic;
	signal Nor258500_o0 : std_logic;
	signal And258520_o0 : std_logic;
	signal Or258540_o0 : std_logic;
	signal Or258560_o0 : std_logic;
	signal Or258580_o0 : std_logic;
	signal And258600_o0 : std_logic;
	signal Or258620_o0 : std_logic;
	signal And258640_o0 : std_logic;
	signal And258660_o0 : std_logic;
	signal Or258680_o0 : std_logic;
	signal And258700_o0 : std_logic;
	signal And258720_o0 : std_logic;
	signal Or258740_o0 : std_logic;
	signal And258760_o0 : std_logic;
	signal And258780_o0 : std_logic;
	signal Or258800_o0 : std_logic;
	signal And258820_o0 : std_logic;
	signal Or258840_o0 : std_logic;
	signal And258860_o0 : std_logic;
	signal And258880_o0 : std_logic;
	signal And258900_o0 : std_logic;
	signal Or258920_o0 : std_logic;
	signal And258940_o0 : std_logic;
	signal And258960_o0 : std_logic;
	signal And258980_o0 : std_logic;
	signal Or259000_o0 : std_logic;
	signal And259020_o0 : std_logic;
	signal And259040_o0 : std_logic;
	signal And259060_o0 : std_logic;
	signal Or259080_o0 : std_logic;
	signal And259100_o0 : std_logic;
	signal Or259120_o0 : std_logic;
	signal And259140_o0 : std_logic;
	signal Or259160_o0 : std_logic;
	signal And259180_o0 : std_logic;
	signal And259200_o0 : std_logic;
	signal Or259220_o0 : std_logic;
	signal And259240_o0 : std_logic;
	signal And259260_o0 : std_logic;
	signal And259280_o0 : std_logic;
	signal And259300_o0 : std_logic;
	signal Or259320_o0 : std_logic;
	signal Or259340_o0 : std_logic;
	signal Or259360_o0 : std_logic;
	signal And259380_o0 : std_logic;
	signal And259400_o0 : std_logic;
	signal And259420_o0 : std_logic;
	signal Or259440_o0 : std_logic;
	signal And259460_o0 : std_logic;
	signal Or259480_o0 : std_logic;
	signal And259500_o0 : std_logic;
	signal And259520_o0 : std_logic;
	signal And259540_o0 : std_logic;
	signal Or259560_o0 : std_logic;
	signal And259580_o0 : std_logic;
	signal Or259600_o0 : std_logic;
	signal And259620_o0 : std_logic;
	signal And259640_o0 : std_logic;
	signal Or259660_o0 : std_logic;
	signal And259680_o0 : std_logic;
	signal And259700_o0 : std_logic;
	signal Or259720_o0 : std_logic;
	signal Or259740_o0 : std_logic;
	signal And259760_o0 : std_logic;
	signal Or259780_o0 : std_logic;
	signal And259800_o0 : std_logic;
	signal And259820_o0 : std_logic;
	signal Or259840_o0 : std_logic;
	signal Or259860_o0 : std_logic;
	signal And259880_o0 : std_logic;
	signal And259900_o0 : std_logic;
	signal And259920_o0 : std_logic;
	signal Or259940_o0 : std_logic;
	signal And259960_o0 : std_logic;
	signal And259980_o0 : std_logic;
	signal Or260000_o0 : std_logic;
	signal And260020_o0 : std_logic;
	signal And260040_o0 : std_logic;
	signal Or260060_o0 : std_logic;
	signal Or260080_o0 : std_logic;
	signal And260100_o0 : std_logic;
	signal And260120_o0 : std_logic;
	signal And260140_o0 : std_logic;
	signal Or260160_o0 : std_logic;
	signal Or260180_o0 : std_logic;
	signal Or260200_o0 : std_logic;
	signal Or260220_o0 : std_logic;
	signal And260240_o0 : std_logic;
	signal Or260260_o0 : std_logic;
	signal And260280_o0 : std_logic;
	signal Or260300_o0 : std_logic;
	signal And260320_o0 : std_logic;
	signal And260340_o0 : std_logic;
	signal Or260360_o0 : std_logic;
	signal And260380_o0 : std_logic;
	signal And260400_o0 : std_logic;
	signal And260420_o0 : std_logic;
	signal Or260440_o0 : std_logic;
	signal And260460_o0 : std_logic;
	signal And260480_o0 : std_logic;
	signal And260500_o0 : std_logic;
	signal And260520_o0 : std_logic;
	signal Or260540_o0 : std_logic;
	signal And260560_o0 : std_logic;
	signal Or260580_o0 : std_logic;
	signal And260600_o0 : std_logic;
	signal And260620_o0 : std_logic;
	signal Or260640_o0 : std_logic;
	signal And260660_o0 : std_logic;
	signal Nor260680_o0 : std_logic;
	signal And260700_o0 : std_logic;
	signal And260720_o0 : std_logic;
	signal Or260740_o0 : std_logic;
	signal And260760_o0 : std_logic;
	signal And260780_o0 : std_logic;
	signal And260800_o0 : std_logic;
	signal Or260820_o0 : std_logic;
	signal And260840_o0 : std_logic;
	signal And260860_o0 : std_logic;
	signal And260880_o0 : std_logic;
	signal And260900_o0 : std_logic;
	signal Or260920_o0 : std_logic;
	signal And260940_o0 : std_logic;
	signal And260960_o0 : std_logic;
	signal And260980_o0 : std_logic;
	signal Or261000_o0 : std_logic;
	signal And261020_o0 : std_logic;
	signal And261040_o0 : std_logic;
	signal Or261060_o0 : std_logic;
	signal And261080_o0 : std_logic;
	signal And261100_o0 : std_logic;
	signal Or261120_o0 : std_logic;
	signal And261140_o0 : std_logic;
	signal And261160_o0 : std_logic;
	signal And261180_o0 : std_logic;
	signal Or261200_o0 : std_logic;
	signal And261220_o0 : std_logic;
	signal And261240_o0 : std_logic;
	signal And261260_o0 : std_logic;
	signal Or261280_o0 : std_logic;
	signal And261300_o0 : std_logic;
	signal And261320_o0 : std_logic;
	signal Or261340_o0 : std_logic;
	signal Or261360_o0 : std_logic;
	signal And261380_o0 : std_logic;
	signal And261400_o0 : std_logic;
	signal And261420_o0 : std_logic;
	signal Or261440_o0 : std_logic;
	signal And261460_o0 : std_logic;
	signal And261480_o0 : std_logic;
	signal And261500_o0 : std_logic;
	signal Or261520_o0 : std_logic;
	signal And261540_o0 : std_logic;
	signal And261560_o0 : std_logic;
	signal Or261580_o0 : std_logic;
	signal And261600_o0 : std_logic;
	signal And261620_o0 : std_logic;
	signal And261640_o0 : std_logic;
	signal And261660_o0 : std_logic;
	signal And261680_o0 : std_logic;
	signal And261700_o0 : std_logic;
	signal And261720_o0 : std_logic;
	signal Or261740_o0 : std_logic;
	signal And261760_o0 : std_logic;
	signal Or261780_o0 : std_logic;
	signal And261800_o0 : std_logic;
	signal And261820_o0 : std_logic;
	signal Or261840_o0 : std_logic;
	signal And261860_o0 : std_logic;
	signal And261880_o0 : std_logic;
	signal Or261900_o0 : std_logic;
	signal And261920_o0 : std_logic;
	signal And261940_o0 : std_logic;
	signal And261960_o0 : std_logic;
	signal And261980_o0 : std_logic;
	signal Or262000_o0 : std_logic;
	signal And262020_o0 : std_logic;
	signal And262040_o0 : std_logic;
	signal And262060_o0 : std_logic;
	signal Or262080_o0 : std_logic;
	signal And262100_o0 : std_logic;
	signal And262120_o0 : std_logic;
	signal Or262140_o0 : std_logic;
	signal And262160_o0 : std_logic;
	signal And262180_o0 : std_logic;
	signal Or262200_o0 : std_logic;
	signal And262220_o0 : std_logic;
	signal And262240_o0 : std_logic;
	signal Or262260_o0 : std_logic;
	signal And262280_o0 : std_logic;
	signal And262300_o0 : std_logic;
	signal Or262320_o0 : std_logic;
	signal And262340_o0 : std_logic;
	signal And262360_o0 : std_logic;
	signal Or262380_o0 : std_logic;
	signal And262400_o0 : std_logic;
	signal And262420_o0 : std_logic;
	signal Nor262440_o0 : std_logic;
	signal And262460_o0 : std_logic;
	signal And262480_o0 : std_logic;
	signal And262500_o0 : std_logic;
	signal Or262520_o0 : std_logic;
	signal And262540_o0 : std_logic;
	signal Or262560_o0 : std_logic;
	signal And262580_o0 : std_logic;
	signal Or262600_o0 : std_logic;
	signal And262620_o0 : std_logic;
	signal Or262640_o0 : std_logic;
	signal Or262660_o0 : std_logic;
	signal And262680_o0 : std_logic;
	signal And262700_o0 : std_logic;
	signal And262720_o0 : std_logic;
	signal And262740_o0 : std_logic;
	signal And262760_o0 : std_logic;
	signal Or262780_o0 : std_logic;
	signal Or262800_o0 : std_logic;
	signal And262820_o0 : std_logic;
	signal And262840_o0 : std_logic;
	signal And262860_o0 : std_logic;
	signal Or262880_o0 : std_logic;
	signal And262900_o0 : std_logic;
	signal And262920_o0 : std_logic;
	signal Or262940_o0 : std_logic;
	signal And262960_o0 : std_logic;
	signal And262980_o0 : std_logic;
	signal And263000_o0 : std_logic;
	signal And263020_o0 : std_logic;
	signal And263040_o0 : std_logic;
	signal Or263060_o0 : std_logic;
	signal And263080_o0 : std_logic;
	signal And263100_o0 : std_logic;
	signal And263120_o0 : std_logic;
	signal Or263140_o0 : std_logic;
	signal And263160_o0 : std_logic;
	signal And263180_o0 : std_logic;
	signal And263200_o0 : std_logic;
	signal And263220_o0 : std_logic;
	signal Or263240_o0 : std_logic;
	signal Nor263260_o0 : std_logic;
	signal And263280_o0 : std_logic;
	signal And263300_o0 : std_logic;
	signal Or263320_o0 : std_logic;
	signal And263340_o0 : std_logic;
	signal And263360_o0 : std_logic;
	signal Or263380_o0 : std_logic;
	signal And263400_o0 : std_logic;
	signal Or263420_o0 : std_logic;
	signal And263440_o0 : std_logic;
	signal And263460_o0 : std_logic;
	signal And263480_o0 : std_logic;
	signal Or263500_o0 : std_logic;
	signal And263520_o0 : std_logic;
	signal Or263540_o0 : std_logic;
	signal And263560_o0 : std_logic;
	signal And263580_o0 : std_logic;
	signal And263600_o0 : std_logic;
	signal Or263620_o0 : std_logic;
	signal And263640_o0 : std_logic;
	signal And263660_o0 : std_logic;
	signal Or263680_o0 : std_logic;
	signal Or263700_o0 : std_logic;
	signal Or263720_o0 : std_logic;
	signal And263740_o0 : std_logic;
	signal Or263760_o0 : std_logic;
	signal And263780_o0 : std_logic;
	signal And263800_o0 : std_logic;
	signal And263820_o0 : std_logic;
	signal Or263840_o0 : std_logic;
	signal And263860_o0 : std_logic;
	signal And263880_o0 : std_logic;
	signal Or263900_o0 : std_logic;
	signal And263920_o0 : std_logic;
	signal Or263940_o0 : std_logic;
	signal And263960_o0 : std_logic;
	signal And263980_o0 : std_logic;
	signal And264000_o0 : std_logic;
	signal And264020_o0 : std_logic;
	signal Or264040_o0 : std_logic;
	signal Or264060_o0 : std_logic;
	signal And264080_o0 : std_logic;
	signal And264100_o0 : std_logic;
	signal And264120_o0 : std_logic;
	signal Or264140_o0 : std_logic;
	signal And264160_o0 : std_logic;
	signal And264180_o0 : std_logic;
	signal And264200_o0 : std_logic;
	signal Or264220_o0 : std_logic;
	signal And264240_o0 : std_logic;
	signal And264260_o0 : std_logic;
	signal And264280_o0 : std_logic;
	signal Or264300_o0 : std_logic;
	signal Or264320_o0 : std_logic;
	signal And264340_o0 : std_logic;
	signal And264360_o0 : std_logic;
	signal Nor264380_o0 : std_logic;
	signal And264400_o0 : std_logic;
	signal Or264420_o0 : std_logic;
	signal And264440_o0 : std_logic;
	signal Or264460_o0 : std_logic;
	signal And264480_o0 : std_logic;
	signal And264500_o0 : std_logic;
	signal And264520_o0 : std_logic;
	signal And264540_o0 : std_logic;
	signal Or264560_o0 : std_logic;
	signal Or264580_o0 : std_logic;
	signal Or264600_o0 : std_logic;
	signal And264620_o0 : std_logic;
	signal And264640_o0 : std_logic;
	signal Or264660_o0 : std_logic;
	signal And264680_o0 : std_logic;
	signal Or264700_o0 : std_logic;
	signal And264720_o0 : std_logic;
	signal And264740_o0 : std_logic;
	signal Or264760_o0 : std_logic;
	signal Or264780_o0 : std_logic;
	signal And264800_o0 : std_logic;
	signal And264820_o0 : std_logic;
	signal Or264840_o0 : std_logic;
	signal Or264860_o0 : std_logic;
	signal Or264880_o0 : std_logic;
	signal And264900_o0 : std_logic;
	signal Or264920_o0 : std_logic;
	signal And264940_o0 : std_logic;
	signal And264960_o0 : std_logic;
	signal And264980_o0 : std_logic;
	signal Or265000_o0 : std_logic;
	signal And265020_o0 : std_logic;
	signal And265040_o0 : std_logic;
	signal And265060_o0 : std_logic;
	signal And265080_o0 : std_logic;
	signal And265100_o0 : std_logic;
	signal And265120_o0 : std_logic;
	signal Or265140_o0 : std_logic;
	signal And265160_o0 : std_logic;
	signal And265180_o0 : std_logic;
	signal And265200_o0 : std_logic;
	signal And265220_o0 : std_logic;
	signal And265240_o0 : std_logic;
	signal And265260_o0 : std_logic;
	signal And265280_o0 : std_logic;
	signal And265300_o0 : std_logic;
	signal And265320_o0 : std_logic;
	signal And265340_o0 : std_logic;
	signal Or265360_o0 : std_logic;
	signal Or265380_o0 : std_logic;
	signal Or265400_o0 : std_logic;
	signal Or265420_o0 : std_logic;
	signal And265440_o0 : std_logic;
	signal And265460_o0 : std_logic;
	signal Or265480_o0 : std_logic;
	signal Or265500_o0 : std_logic;
	signal And265520_o0 : std_logic;
	signal And265540_o0 : std_logic;
	signal Or265560_o0 : std_logic;
	signal And265580_o0 : std_logic;
	signal And265600_o0 : std_logic;
	signal Or265620_o0 : std_logic;
	signal And265640_o0 : std_logic;
	signal And265660_o0 : std_logic;
	signal And265680_o0 : std_logic;
	signal And265700_o0 : std_logic;
	signal And265720_o0 : std_logic;
	signal And265740_o0 : std_logic;
	signal Or265760_o0 : std_logic;
	signal And265780_o0 : std_logic;
	signal And265800_o0 : std_logic;
	signal Or265820_o0 : std_logic;
	signal And265840_o0 : std_logic;
	signal And265860_o0 : std_logic;
	signal Or265880_o0 : std_logic;
	signal And265900_o0 : std_logic;
	signal And265920_o0 : std_logic;
	signal Or265940_o0 : std_logic;
	signal And265960_o0 : std_logic;
	signal And265980_o0 : std_logic;
	signal And266000_o0 : std_logic;
	signal And266020_o0 : std_logic;
	signal Or266040_o0 : std_logic;
	signal And266060_o0 : std_logic;
	signal Or266080_o0 : std_logic;
	signal And266100_o0 : std_logic;
	signal And266120_o0 : std_logic;
	signal Or266140_o0 : std_logic;
	signal And266160_o0 : std_logic;
	signal And266180_o0 : std_logic;
	signal And266200_o0 : std_logic;
	signal Or266220_o0 : std_logic;
	signal And266240_o0 : std_logic;
	signal And266260_o0 : std_logic;
	signal And266280_o0 : std_logic;
	signal Or266300_o0 : std_logic;
	signal And266320_o0 : std_logic;
	signal And266340_o0 : std_logic;
	signal Or266360_o0 : std_logic;
	signal And266380_o0 : std_logic;
	signal And266400_o0 : std_logic;
	signal And266420_o0 : std_logic;
	signal And266440_o0 : std_logic;
	signal Or266460_o0 : std_logic;
	signal And266480_o0 : std_logic;
	signal Or266500_o0 : std_logic;
	signal And266520_o0 : std_logic;
	signal Or266540_o0 : std_logic;
	signal And266560_o0 : std_logic;
	signal Nor266580_o0 : std_logic;
	signal Or266600_o0 : std_logic;
	signal And266620_o0 : std_logic;
	signal Or266640_o0 : std_logic;
	signal And266660_o0 : std_logic;
	signal And266680_o0 : std_logic;
	signal Or266700_o0 : std_logic;
	signal And266720_o0 : std_logic;
	signal Or266740_o0 : std_logic;
	signal And266760_o0 : std_logic;
	signal Or266780_o0 : std_logic;
	signal And266800_o0 : std_logic;
	signal And266820_o0 : std_logic;
	signal And266840_o0 : std_logic;
	signal Or266860_o0 : std_logic;
	signal And266880_o0 : std_logic;
	signal Or266900_o0 : std_logic;
	signal And266920_o0 : std_logic;
	signal Or266940_o0 : std_logic;
	signal Or266960_o0 : std_logic;
	signal And266980_o0 : std_logic;
	signal And267000_o0 : std_logic;
	signal And267020_o0 : std_logic;
	signal And267040_o0 : std_logic;
	signal Or267060_o0 : std_logic;
	signal And267080_o0 : std_logic;
	signal And267100_o0 : std_logic;
	signal And267120_o0 : std_logic;
	signal And267140_o0 : std_logic;
	signal Or267160_o0 : std_logic;
	signal And267180_o0 : std_logic;
	signal And267200_o0 : std_logic;
	signal And267220_o0 : std_logic;
	signal Or267240_o0 : std_logic;
	signal And267260_o0 : std_logic;
	signal Or267280_o0 : std_logic;
	signal And267300_o0 : std_logic;
	signal And267320_o0 : std_logic;
	signal Or267340_o0 : std_logic;
	signal And267360_o0 : std_logic;
	signal And267380_o0 : std_logic;
	signal Or267400_o0 : std_logic;
	signal And267420_o0 : std_logic;
	signal And267440_o0 : std_logic;
	signal And267460_o0 : std_logic;
	signal Or267480_o0 : std_logic;
	signal And267500_o0 : std_logic;
	signal And267520_o0 : std_logic;
	signal And267540_o0 : std_logic;
	signal And267560_o0 : std_logic;
	signal Or267580_o0 : std_logic;
	signal And267600_o0 : std_logic;
	signal Nor267620_o0 : std_logic;
	signal And267640_o0 : std_logic;
	signal Or267660_o0 : std_logic;
	signal And267680_o0 : std_logic;
	signal And267700_o0 : std_logic;
	signal And267720_o0 : std_logic;
	signal Or267740_o0 : std_logic;
	signal And267760_o0 : std_logic;
	signal And267780_o0 : std_logic;
	signal And267800_o0 : std_logic;
	signal Or267820_o0 : std_logic;
	signal And267840_o0 : std_logic;
	signal And267860_o0 : std_logic;
	signal And267880_o0 : std_logic;
	signal Or267900_o0 : std_logic;
	signal And267920_o0 : std_logic;
	signal Or267940_o0 : std_logic;
	signal And267960_o0 : std_logic;
	signal Or267980_o0 : std_logic;
	signal And268000_o0 : std_logic;
	signal And268020_o0 : std_logic;
	signal Or268040_o0 : std_logic;
	signal And268060_o0 : std_logic;
	signal Or268080_o0 : std_logic;
	signal And268100_o0 : std_logic;
	signal And268120_o0 : std_logic;
	signal Or268140_o0 : std_logic;
	signal Or268160_o0 : std_logic;
	signal And268180_o0 : std_logic;
	signal And268200_o0 : std_logic;
	signal And268220_o0 : std_logic;
	signal Or268240_o0 : std_logic;
	signal And268260_o0 : std_logic;
	signal And268280_o0 : std_logic;
	signal Or268300_o0 : std_logic;
	signal And268320_o0 : std_logic;
	signal And268340_o0 : std_logic;
	signal Or268360_o0 : std_logic;
	signal And268380_o0 : std_logic;
	signal And268400_o0 : std_logic;
	signal Or268420_o0 : std_logic;
	signal And268440_o0 : std_logic;
	signal And268460_o0 : std_logic;
	signal And268480_o0 : std_logic;
	signal And268500_o0 : std_logic;
	signal Or268520_o0 : std_logic;
	signal And268540_o0 : std_logic;
	signal And268560_o0 : std_logic;
	signal And268580_o0 : std_logic;
	signal Or268600_o0 : std_logic;
	signal And268620_o0 : std_logic;
	signal And268640_o0 : std_logic;
	signal And268660_o0 : std_logic;
	signal And268680_o0 : std_logic;
	signal And268700_o0 : std_logic;
	signal And268720_o0 : std_logic;
	signal Or268740_o0 : std_logic;
	signal And268760_o0 : std_logic;
	signal And268780_o0 : std_logic;
	signal And268800_o0 : std_logic;
	signal Or268820_o0 : std_logic;
	signal And268840_o0 : std_logic;
	signal And268860_o0 : std_logic;
	signal And268880_o0 : std_logic;
	signal Or268900_o0 : std_logic;
	signal And268920_o0 : std_logic;
	signal And268940_o0 : std_logic;
	signal And268960_o0 : std_logic;
	signal And268980_o0 : std_logic;
	signal Or269000_o0 : std_logic;
	signal And269020_o0 : std_logic;
	signal And269040_o0 : std_logic;
	signal Or269060_o0 : std_logic;
	signal And269080_o0 : std_logic;
	signal And269100_o0 : std_logic;
	signal Or269120_o0 : std_logic;
	signal And269140_o0 : std_logic;
	signal And269160_o0 : std_logic;
	signal Or269180_o0 : std_logic;
	signal And269200_o0 : std_logic;
	signal Nor269220_o0 : std_logic;
	signal And269240_o0 : std_logic;
	signal And269260_o0 : std_logic;
	signal And269280_o0 : std_logic;
	signal Or269300_o0 : std_logic;
	signal And269320_o0 : std_logic;
	signal Xor269340_o0 : std_logic;
	signal And269360_o0 : std_logic;
	signal And269380_o0 : std_logic;
	signal And269400_o0 : std_logic;
	signal And269420_o0 : std_logic;
	signal Or269440_o0 : std_logic;
	signal And269460_o0 : std_logic;
	signal Nor269480_o0 : std_logic;
	signal And269500_o0 : std_logic;
	signal Or269520_o0 : std_logic;
	signal And269540_o0 : std_logic;
	signal And269560_o0 : std_logic;
	signal And269580_o0 : std_logic;
	signal And269600_o0 : std_logic;
	signal And269620_o0 : std_logic;
	signal Or269640_o0 : std_logic;
	signal And269660_o0 : std_logic;
	signal And269680_o0 : std_logic;
	signal And269700_o0 : std_logic;
	signal And269720_o0 : std_logic;
	signal And269740_o0 : std_logic;
	signal And269760_o0 : std_logic;
	signal And269780_o0 : std_logic;
	signal Or269800_o0 : std_logic;
	signal And269820_o0 : std_logic;
	signal And269840_o0 : std_logic;
	signal And269860_o0 : std_logic;
	signal And269880_o0 : std_logic;
	signal Or269900_o0 : std_logic;
	signal And269920_o0 : std_logic;
	signal And269940_o0 : std_logic;
	signal And269960_o0 : std_logic;
	signal Or269980_o0 : std_logic;
	signal And270000_o0 : std_logic;
	signal And270020_o0 : std_logic;
	signal Or270040_o0 : std_logic;
	signal And270060_o0 : std_logic;
	signal And270080_o0 : std_logic;
	signal And270100_o0 : std_logic;
	signal And270120_o0 : std_logic;
	signal Or270140_o0 : std_logic;
	signal And270160_o0 : std_logic;
	signal And270180_o0 : std_logic;
	signal And270200_o0 : std_logic;
	signal Or270220_o0 : std_logic;
	signal And270240_o0 : std_logic;
	signal And270260_o0 : std_logic;
	signal Or270280_o0 : std_logic;
	signal And270300_o0 : std_logic;
	signal Or270320_o0 : std_logic;
	signal And270340_o0 : std_logic;
	signal And270360_o0 : std_logic;
	signal Or270380_o0 : std_logic;
	signal And270400_o0 : std_logic;
	signal And270420_o0 : std_logic;
	signal And270440_o0 : std_logic;
	signal And270460_o0 : std_logic;
	signal Or270480_o0 : std_logic;
	signal And270500_o0 : std_logic;
	signal And270520_o0 : std_logic;
	signal And270540_o0 : std_logic;
	signal And270560_o0 : std_logic;
	signal And270580_o0 : std_logic;
	signal Or270600_o0 : std_logic;
	signal And270620_o0 : std_logic;
	signal And270640_o0 : std_logic;
	signal And270660_o0 : std_logic;
	signal Or270680_o0 : std_logic;
	signal And270700_o0 : std_logic;
	signal And270720_o0 : std_logic;
	signal Or270740_o0 : std_logic;
	signal And270760_o0 : std_logic;
	signal And270780_o0 : std_logic;
	signal And270800_o0 : std_logic;
	signal Or270820_o0 : std_logic;
	signal And270840_o0 : std_logic;
	signal Or270860_o0 : std_logic;
	signal Or270880_o0 : std_logic;
	signal And270900_o0 : std_logic;
	signal And270920_o0 : std_logic;
	signal Or270940_o0 : std_logic;
	signal And270960_o0 : std_logic;
	signal And270980_o0 : std_logic;
	signal And271000_o0 : std_logic;
	signal And271020_o0 : std_logic;
	signal Or271040_o0 : std_logic;
	signal And271060_o0 : std_logic;
	signal And271080_o0 : std_logic;
	signal And271100_o0 : std_logic;
	signal And271120_o0 : std_logic;
	signal Or271140_o0 : std_logic;
	signal And271160_o0 : std_logic;
	signal And271180_o0 : std_logic;
	signal And271200_o0 : std_logic;
	signal And271220_o0 : std_logic;
	signal Or271240_o0 : std_logic;
	signal And271260_o0 : std_logic;
	signal And271280_o0 : std_logic;
	signal Or271300_o0 : std_logic;
	signal And271320_o0 : std_logic;
	signal Or271340_o0 : std_logic;
	signal And271360_o0 : std_logic;
	signal And271380_o0 : std_logic;
	signal And271400_o0 : std_logic;
	signal And271420_o0 : std_logic;
	signal And271440_o0 : std_logic;
	signal And271460_o0 : std_logic;
	signal And271480_o0 : std_logic;
	signal Or271500_o0 : std_logic;
	signal And271520_o0 : std_logic;
	signal Or271540_o0 : std_logic;
	signal And271560_o0 : std_logic;
	signal And271580_o0 : std_logic;
	signal And271600_o0 : std_logic;
	signal Or271620_o0 : std_logic;
	signal And271640_o0 : std_logic;
	signal And271660_o0 : std_logic;
	signal And271680_o0 : std_logic;
	signal And271700_o0 : std_logic;
	signal And271720_o0 : std_logic;
	signal And271740_o0 : std_logic;
	signal Or271760_o0 : std_logic;
	signal And271780_o0 : std_logic;
	signal And271800_o0 : std_logic;
	signal And271820_o0 : std_logic;
	signal Or271840_o0 : std_logic;
	signal And271860_o0 : std_logic;
	signal Or271880_o0 : std_logic;
	signal And271900_o0 : std_logic;
	signal Or271920_o0 : std_logic;
	signal And271940_o0 : std_logic;
	signal And271960_o0 : std_logic;
	signal Or271980_o0 : std_logic;
	signal And272000_o0 : std_logic;
	signal And272020_o0 : std_logic;
	signal And272040_o0 : std_logic;
	signal Or272060_o0 : std_logic;
	signal And272080_o0 : std_logic;
	signal And272100_o0 : std_logic;
	signal And272120_o0 : std_logic;
	signal Or272140_o0 : std_logic;
	signal And272160_o0 : std_logic;
	signal And272180_o0 : std_logic;
	signal And272200_o0 : std_logic;
	signal And272220_o0 : std_logic;
	signal And272240_o0 : std_logic;
	signal And272260_o0 : std_logic;
	signal Or272280_o0 : std_logic;
	signal Nor272300_o0 : std_logic;
	signal And272320_o0 : std_logic;
	signal And272340_o0 : std_logic;
	signal And272360_o0 : std_logic;
	signal And272380_o0 : std_logic;
	signal And272400_o0 : std_logic;
	signal Or272420_o0 : std_logic;
	signal And272440_o0 : std_logic;
	signal And272460_o0 : std_logic;
	signal And272480_o0 : std_logic;
	signal Nor272500_o0 : std_logic;
	signal And272520_o0 : std_logic;
	signal And272540_o0 : std_logic;
	signal And272560_o0 : std_logic;
	signal And272580_o0 : std_logic;
	signal And272600_o0 : std_logic;
	signal And272620_o0 : std_logic;
	signal And272640_o0 : std_logic;
	signal And272660_o0 : std_logic;
	signal Or272680_o0 : std_logic;
	signal And272700_o0 : std_logic;
	signal And272720_o0 : std_logic;
	signal Or272740_o0 : std_logic;
	signal And272760_o0 : std_logic;
	signal Or272780_o0 : std_logic;
	signal And272800_o0 : std_logic;
	signal And272820_o0 : std_logic;
	signal And272840_o0 : std_logic;
	signal Nor272860_o0 : std_logic;
	signal And272880_o0 : std_logic;
	signal Or272900_o0 : std_logic;
	signal Or272920_o0 : std_logic;
	signal And272940_o0 : std_logic;
	signal And272960_o0 : std_logic;
	signal And272980_o0 : std_logic;
	signal And273000_o0 : std_logic;
	signal And273020_o0 : std_logic;
	signal Or273040_o0 : std_logic;
	signal And273060_o0 : std_logic;
	signal And273080_o0 : std_logic;
	signal Or273100_o0 : std_logic;
	signal Or273120_o0 : std_logic;
	signal Or273140_o0 : std_logic;
	signal And273160_o0 : std_logic;
	signal And273180_o0 : std_logic;
	signal And273200_o0 : std_logic;
	signal Or273220_o0 : std_logic;
	signal And273240_o0 : std_logic;
	signal And273260_o0 : std_logic;
	signal Or273280_o0 : std_logic;
	signal And273300_o0 : std_logic;
	signal And273320_o0 : std_logic;
	signal And273340_o0 : std_logic;
	signal And273360_o0 : std_logic;
	signal Or273380_o0 : std_logic;
	signal And273400_o0 : std_logic;
	signal Or273420_o0 : std_logic;
	signal And273440_o0 : std_logic;
	signal And273460_o0 : std_logic;
	signal Or273480_o0 : std_logic;
	signal And273500_o0 : std_logic;
	signal And273520_o0 : std_logic;
	signal And273540_o0 : std_logic;
	signal Or273560_o0 : std_logic;
	signal And273580_o0 : std_logic;
	signal And273600_o0 : std_logic;
	signal And273620_o0 : std_logic;
	signal Or273640_o0 : std_logic;
	signal And273660_o0 : std_logic;
	signal And273680_o0 : std_logic;
	signal Or273700_o0 : std_logic;
	signal And273720_o0 : std_logic;
	signal And273740_o0 : std_logic;
	signal Nor273760_o0 : std_logic;
	signal And273780_o0 : std_logic;
	signal And273800_o0 : std_logic;
	signal Or273820_o0 : std_logic;
	signal And273840_o0 : std_logic;
	signal And273860_o0 : std_logic;
	signal And273880_o0 : std_logic;
	signal And273900_o0 : std_logic;
	signal Or273920_o0 : std_logic;
	signal And273940_o0 : std_logic;
	signal And273960_o0 : std_logic;
	signal Nor273980_o0 : std_logic;
	signal Nor274000_o0 : std_logic;
	signal And274020_o0 : std_logic;
	signal And274040_o0 : std_logic;
	signal And274060_o0 : std_logic;
	signal And274080_o0 : std_logic;
	signal And274100_o0 : std_logic;
	signal And274120_o0 : std_logic;
	signal And274140_o0 : std_logic;
	signal And274160_o0 : std_logic;
	signal Or274180_o0 : std_logic;
	signal And274200_o0 : std_logic;
	signal And274220_o0 : std_logic;
	signal And274240_o0 : std_logic;
	signal And274260_o0 : std_logic;
	signal Or274280_o0 : std_logic;
	signal And274300_o0 : std_logic;
	signal And274320_o0 : std_logic;
	signal And274340_o0 : std_logic;
	signal Or274360_o0 : std_logic;
	signal And274380_o0 : std_logic;
	signal And274400_o0 : std_logic;
	signal Or274420_o0 : std_logic;
	signal And274440_o0 : std_logic;
	signal Or274460_o0 : std_logic;
	signal And274480_o0 : std_logic;
	signal And274500_o0 : std_logic;
	signal And274520_o0 : std_logic;
	signal Or274540_o0 : std_logic;
	signal Or274560_o0 : std_logic;
	signal Or274580_o0 : std_logic;
	signal And274600_o0 : std_logic;
	signal And274620_o0 : std_logic;
	signal And274640_o0 : std_logic;
	signal And274660_o0 : std_logic;
	signal Or274680_o0 : std_logic;
	signal And274700_o0 : std_logic;
	signal Or274720_o0 : std_logic;
	signal And274740_o0 : std_logic;
	signal Or274760_o0 : std_logic;
	signal And274780_o0 : std_logic;
	signal And274800_o0 : std_logic;
	signal And274820_o0 : std_logic;
	signal And274840_o0 : std_logic;
	signal And274860_o0 : std_logic;
	signal And274880_o0 : std_logic;
	signal Or274900_o0 : std_logic;
	signal And274920_o0 : std_logic;
	signal Xor274940_o0 : std_logic;
	signal And274960_o0 : std_logic;
	signal And274980_o0 : std_logic;
	signal And275000_o0 : std_logic;
	signal Or275020_o0 : std_logic;
	signal Or275040_o0 : std_logic;
	signal And275060_o0 : std_logic;
	signal And275080_o0 : std_logic;
	signal Or275100_o0 : std_logic;
	signal And275120_o0 : std_logic;
	signal Or275140_o0 : std_logic;
	signal And275160_o0 : std_logic;
	signal And275180_o0 : std_logic;
	signal Or275200_o0 : std_logic;
	signal And275220_o0 : std_logic;
	signal And275240_o0 : std_logic;
	signal And275260_o0 : std_logic;
	signal Or275280_o0 : std_logic;
	signal And275300_o0 : std_logic;
	signal Or275320_o0 : std_logic;
	signal And275340_o0 : std_logic;
	signal And275360_o0 : std_logic;
	signal And275380_o0 : std_logic;
	signal Or275400_o0 : std_logic;
	signal And275420_o0 : std_logic;
	signal And275440_o0 : std_logic;
	signal And275460_o0 : std_logic;
	signal And275480_o0 : std_logic;
	signal Or275500_o0 : std_logic;
	signal And275520_o0 : std_logic;
	signal And275540_o0 : std_logic;
	signal And275560_o0 : std_logic;
	signal And275580_o0 : std_logic;
	signal Or275600_o0 : std_logic;
	signal And275620_o0 : std_logic;
	signal And275640_o0 : std_logic;
	signal And275660_o0 : std_logic;
	signal And275680_o0 : std_logic;
	signal And275700_o0 : std_logic;
	signal And275720_o0 : std_logic;
	signal Nor275740_o0 : std_logic;
	signal And275760_o0 : std_logic;
	signal Or275780_o0 : std_logic;
	signal And275800_o0 : std_logic;
	signal And275820_o0 : std_logic;
	signal Or275840_o0 : std_logic;
	signal And275860_o0 : std_logic;
	signal And275880_o0 : std_logic;
	signal And275900_o0 : std_logic;
	signal Or275920_o0 : std_logic;
	signal And275940_o0 : std_logic;
	signal And275960_o0 : std_logic;
	signal And275980_o0 : std_logic;
	signal And276000_o0 : std_logic;
	signal Or276020_o0 : std_logic;
	signal And276040_o0 : std_logic;
	signal And276060_o0 : std_logic;
	signal And276080_o0 : std_logic;
	signal Or276100_o0 : std_logic;
	signal And276120_o0 : std_logic;
	signal And276140_o0 : std_logic;
	signal Or276160_o0 : std_logic;
	signal And276180_o0 : std_logic;
	signal Or276200_o0 : std_logic;
	signal And276220_o0 : std_logic;
	signal And276240_o0 : std_logic;
	signal And276260_o0 : std_logic;
	signal Or276280_o0 : std_logic;
	signal And276300_o0 : std_logic;
	signal And276320_o0 : std_logic;
	signal And276340_o0 : std_logic;
	signal And276360_o0 : std_logic;
	signal And276380_o0 : std_logic;
	signal And276400_o0 : std_logic;
	signal And276420_o0 : std_logic;
	signal Or276440_o0 : std_logic;
	signal And276460_o0 : std_logic;
	signal And276480_o0 : std_logic;
	signal Or276500_o0 : std_logic;
	signal And276520_o0 : std_logic;
	signal And276540_o0 : std_logic;
	signal And276560_o0 : std_logic;
	signal And276580_o0 : std_logic;
	signal Or276600_o0 : std_logic;
	signal And276620_o0 : std_logic;
	signal And276640_o0 : std_logic;
	signal And276660_o0 : std_logic;
	signal And276680_o0 : std_logic;
	signal Or276700_o0 : std_logic;
	signal And276720_o0 : std_logic;
	signal And276740_o0 : std_logic;
	signal And276760_o0 : std_logic;
	signal And276780_o0 : std_logic;
	signal Or276800_o0 : std_logic;
	signal And276820_o0 : std_logic;
	signal And276840_o0 : std_logic;
	signal And276860_o0 : std_logic;
	signal Or276880_o0 : std_logic;
	signal And276900_o0 : std_logic;
	signal And276920_o0 : std_logic;
	signal And276940_o0 : std_logic;
	signal Or276960_o0 : std_logic;
	signal And276980_o0 : std_logic;
	signal And277000_o0 : std_logic;
	signal And277020_o0 : std_logic;
	signal And277040_o0 : std_logic;
	signal Or277060_o0 : std_logic;
	signal And277080_o0 : std_logic;
	signal And277100_o0 : std_logic;
	signal And277120_o0 : std_logic;
	signal And277140_o0 : std_logic;
	signal And277160_o0 : std_logic;
	signal And277180_o0 : std_logic;
	signal And277200_o0 : std_logic;
	signal Or277220_o0 : std_logic;
	signal And277240_o0 : std_logic;
	signal And277260_o0 : std_logic;
	signal And277280_o0 : std_logic;
	signal And277300_o0 : std_logic;
	signal And277320_o0 : std_logic;
	signal Or277340_o0 : std_logic;
	signal And277360_o0 : std_logic;
	signal Or277380_o0 : std_logic;
	signal And277400_o0 : std_logic;
	signal And277420_o0 : std_logic;
	signal And277440_o0 : std_logic;
	signal Or277460_o0 : std_logic;
	signal And277480_o0 : std_logic;
	signal Or277500_o0 : std_logic;
	signal And277520_o0 : std_logic;
	signal Or277540_o0 : std_logic;
	signal And277560_o0 : std_logic;
	signal Or277580_o0 : std_logic;
	signal And277600_o0 : std_logic;
	signal And277620_o0 : std_logic;
	signal And277640_o0 : std_logic;
	signal And277660_o0 : std_logic;
	signal And277680_o0 : std_logic;
	signal Or277700_o0 : std_logic;
	signal And277720_o0 : std_logic;
	signal And277740_o0 : std_logic;
	signal And277760_o0 : std_logic;
	signal Or277780_o0 : std_logic;
	signal And277800_o0 : std_logic;
	signal And277820_o0 : std_logic;
	signal And277840_o0 : std_logic;
	signal And277860_o0 : std_logic;
	signal Or277880_o0 : std_logic;
	signal And277900_o0 : std_logic;
	signal And277920_o0 : std_logic;
	signal Or277940_o0 : std_logic;
	signal And277960_o0 : std_logic;
	signal And277980_o0 : std_logic;
	signal And278000_o0 : std_logic;
	signal Or278020_o0 : std_logic;
	signal And278040_o0 : std_logic;
	signal Or278060_o0 : std_logic;
	signal And278080_o0 : std_logic;
	signal Or279120_o0 : std_logic;
	signal Nor279140_o0 : std_logic;
	signal Nor279160_o0 : std_logic;
	signal And279180_o0 : std_logic;
begin
	----------------------------------
	-- Components interconnect 
	----------------------------------
	Not60 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i0,
			o0 => Not60_o0
		);
		Not80 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			o0 => Not80_o0
		);
		Not100 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i1,
			o0 => Not100_o0
		);
		Not120 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i2,
			o0 => Not120_o0
		);
		Not140 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i3,
			o0 => Not140_o0
		);
		Not160 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			o0 => Not160_o0
		);
		Not180 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			o0 => Not180_o0
		);
		Xor2200 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i15,
			o0 => Xor2200_o0
		);
		Nor2220 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i17,
			o0 => Nor2220_o0
		);
		And2240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i18,
			o0 => And2240_o0
		);
		And2260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2240_o0,
			i1 => i17,
			o0 => And2260_o0
		);
		Or2280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2260_o0,
			i1 => Nor2220_o0,
			o0 => Or2280_o0
		);
		And2300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2280_o0,
			i1 => Xor2200_o0,
			o0 => And2300_o0
		);
		And2320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => i16,
			o0 => And2320_o0
		);
		And2340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2320_o0,
			i1 => i15,
			o0 => And2340_o0
		);
		Or2360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2340_o0,
			i1 => And2300_o0,
			o0 => Or2360_o0
		);
		And2380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2360_o0,
			i1 => Not180_o0,
			o0 => And2380_o0
		);
		And2400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i28,
			i1 => i25,
			o0 => And2400_o0
		);
		And2420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2400_o0,
			i1 => i24,
			o0 => And2420_o0
		);
		Nor2440 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i31,
			i1 => i28,
			o0 => Nor2440_o0
		);
		Or2460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2440_o0,
			i1 => And2420_o0,
			o0 => Or2460_o0
		);
		Or2480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or2460_o0,
			i1 => i15,
			o0 => Or2480_o0
		);
		And2500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2480_o0,
			i1 => i12,
			o0 => And2500_o0
		);
		Or2520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2500_o0,
			i1 => And2380_o0,
			o0 => Or2520_o0
		);
		Not540 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			o0 => Not540_o0
		);
		And2560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not540_o0,
			o0 => And2560_o0
		);
		And2580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => Or2520_o0,
			o0 => And2580_o0
		);
		And2600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => i15,
			o0 => And2600_o0
		);
		Not620 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			o0 => Not620_o0
		);
		And2640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not620_o0,
			o0 => And2640_o0
		);
		And2660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2260_o0,
			i1 => And2640_o0,
			o0 => And2660_o0
		);
		Or2680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2660_o0,
			i1 => And2600_o0,
			o0 => Or2680_o0
		);
		And2700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2680_o0,
			i1 => Not180_o0,
			o0 => And2700_o0
		);
		And2720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2700_o0,
			i1 => i5,
			o0 => And2720_o0
		);
		Or2740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2720_o0,
			i1 => And2580_o0,
			o0 => Or2740_o0
		);
		And2760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2740_o0,
			i1 => Not160_o0,
			o0 => And2760_o0
		);
		And2780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2700_o0,
			i1 => i4,
			o0 => And2780_o0
		);
		Or2800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2780_o0,
			i1 => And2760_o0,
			o0 => Or2800_o0
		);
		And2820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2800_o0,
			i1 => Not140_o0,
			o0 => And2820_o0
		);
		And2840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2700_o0,
			i1 => i3,
			o0 => And2840_o0
		);
		Or2860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2840_o0,
			i1 => And2820_o0,
			o0 => Or2860_o0
		);
		And2880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2860_o0,
			i1 => Not120_o0,
			o0 => And2880_o0
		);
		And2900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2700_o0,
			i1 => i2,
			o0 => And2900_o0
		);
		Or2920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And2900_o0,
			i1 => And2880_o0,
			o0 => Or2920_o0
		);
		And2940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or2920_o0,
			i1 => Not100_o0,
			o0 => And2940_o0
		);
		Xor2960 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i16,
			o0 => Xor2960_o0
		);
		And2980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor2960_o0,
			i1 => Nor2220_o0,
			o0 => And2980_o0
		);
		And21000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2980_o0,
			i1 => i15,
			o0 => And21000_o0
		);
		Or21020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21000_o0,
			i1 => And2660_o0,
			o0 => Or21020_o0
		);
		Not1040 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			o0 => Not1040_o0
		);
		And21060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i16,
			o0 => And21060_o0
		);
		Not1080 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			o0 => Not1080_o0
		);
		And21100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not1080_o0,
			o0 => And21100_o0
		);
		And21120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => And21060_o0,
			o0 => And21120_o0
		);
		Nor21140 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i3,
			i1 => i2,
			o0 => Nor21140_o0
		);
		And21160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not160_o0,
			o0 => And21160_o0
		);
		And21180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21160_o0,
			i1 => Nor21140_o0,
			o0 => And21180_o0
		);
		And21200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21180_o0,
			i1 => And21120_o0,
			o0 => And21200_o0
		);
		Nor21220 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i18,
			o0 => Nor21220_o0
		);
		And21240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => Not1040_o0,
			o0 => And21240_o0
		);
		Nor21260 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i4,
			o0 => Nor21260_o0
		);
		Not1280 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			o0 => Not1280_o0
		);
		And21300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1280_o0,
			i1 => i15,
			o0 => And21300_o0
		);
		And21320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21140_o0,
			i1 => And21300_o0,
			o0 => And21320_o0
		);
		And21340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21320_o0,
			i1 => Nor21260_o0,
			o0 => And21340_o0
		);
		And21360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21340_o0,
			i1 => And21240_o0,
			o0 => And21360_o0
		);
		Or21380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21360_o0,
			i1 => And21200_o0,
			o0 => Or21380_o0
		);
		Or21400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or21380_o0,
			i1 => Or21020_o0,
			o0 => Or21400_o0
		);
		And21420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not180_o0,
			i1 => i1,
			o0 => And21420_o0
		);
		And21440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21420_o0,
			i1 => Or21400_o0,
			o0 => And21440_o0
		);
		Or21460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21440_o0,
			i1 => And2940_o0,
			o0 => Or21460_o0
		);
		And21480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21460_o0,
			i1 => i13,
			o0 => And21480_o0
		);
		Not1500 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			o0 => Not1500_o0
		);
		And21520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1500_o0,
			i1 => i17,
			o0 => And21520_o0
		);
		And21540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21520_o0,
			i1 => i15,
			o0 => And21540_o0
		);
		Xor21560 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not620_o0,
			o0 => Xor21560_o0
		);
		Or21580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Xor21560_o0,
			i1 => And21540_o0,
			o0 => Or21580_o0
		);
		And21600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21580_o0,
			i1 => Not1080_o0,
			o0 => And21600_o0
		);
		Xor21620 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i15,
			o0 => Xor21620_o0
		);
		And21640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i17,
			o0 => And21640_o0
		);
		And21660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => Xor21620_o0,
			o0 => And21660_o0
		);
		Or21680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21660_o0,
			i1 => And21600_o0,
			o0 => Or21680_o0
		);
		And21700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21680_o0,
			i1 => Not1280_o0,
			o0 => And21700_o0
		);
		Or21720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i18,
			o0 => Or21720_o0
		);
		And21740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => i17,
			o0 => And21740_o0
		);
		And21760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21740_o0,
			i1 => Or21720_o0,
			o0 => And21760_o0
		);
		Or21780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21760_o0,
			i1 => And21700_o0,
			o0 => Or21780_o0
		);
		And21800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21780_o0,
			i1 => And2560_o0,
			o0 => And21800_o0
		);
		And21820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => i17,
			o0 => And21820_o0
		);
		Nor21840 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i15,
			o0 => Nor21840_o0
		);
		And21860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => i5,
			o0 => And21860_o0
		);
		And21880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21860_o0,
			i1 => And21820_o0,
			o0 => And21880_o0
		);
		Or21900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21880_o0,
			i1 => And21800_o0,
			o0 => Or21900_o0
		);
		And21920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21900_o0,
			i1 => Not140_o0,
			o0 => And21920_o0
		);
		And21940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not1280_o0,
			o0 => And21940_o0
		);
		And21960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => Nor21220_o0,
			o0 => And21960_o0
		);
		Nor21980 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i5,
			o0 => Nor21980_o0
		);
		And22000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21980_o0,
			i1 => i3,
			o0 => And22000_o0
		);
		And22020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22000_o0,
			i1 => And21960_o0,
			o0 => And22020_o0
		);
		Or22040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22020_o0,
			i1 => And21920_o0,
			o0 => Or22040_o0
		);
		Nor22060 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i2,
			i1 => i1,
			o0 => Nor22060_o0
		);
		Not2080 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			o0 => Not2080_o0
		);
		And22100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => Not160_o0,
			o0 => And22100_o0
		);
		And22120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22100_o0,
			i1 => Not2080_o0,
			o0 => And22120_o0
		);
		And22140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22120_o0,
			i1 => Nor22060_o0,
			o0 => And22140_o0
		);
		And22160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22140_o0,
			i1 => Or22040_o0,
			o0 => And22160_o0
		);
		Or22180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22160_o0,
			i1 => And21480_o0,
			o0 => Or22180_o0
		);
		And22200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22180_o0,
			i1 => Not80_o0,
			o0 => And22200_o0
		);
		And22220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i15,
			o0 => And22220_o0
		);
		And22240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => Not620_o0,
			o0 => And22240_o0
		);
		Or22260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22240_o0,
			i1 => And22220_o0,
			o0 => Or22260_o0
		);
		And22280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22260_o0,
			i1 => Not1040_o0,
			o0 => And22280_o0
		);
		And22300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not620_o0,
			o0 => And22300_o0
		);
		And22320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22300_o0,
			i1 => And2240_o0,
			o0 => And22320_o0
		);
		Or22340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22320_o0,
			i1 => And22280_o0,
			o0 => Or22340_o0
		);
		And22360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22340_o0,
			i1 => Not1280_o0,
			o0 => And22360_o0
		);
		And22380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21720_o0,
			i1 => Not1040_o0,
			o0 => And22380_o0
		);
		And22400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i15,
			o0 => And22400_o0
		);
		And22420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22400_o0,
			i1 => And22380_o0,
			o0 => And22420_o0
		);
		Or22440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22420_o0,
			i1 => And22360_o0,
			o0 => Or22440_o0
		);
		And22460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22440_o0,
			i1 => i13,
			o0 => And22460_o0
		);
		And22480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i13,
			o0 => And22480_o0
		);
		And22500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22480_o0,
			i1 => And21240_o0,
			o0 => And22500_o0
		);
		Or22520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22500_o0,
			i1 => Not2080_o0,
			o0 => Or22520_o0
		);
		Or22540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or22520_o0,
			i1 => And22460_o0,
			o0 => Or22540_o0
		);
		And22560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i12,
			o0 => And22560_o0
		);
		And22580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22560_o0,
			i1 => And2560_o0,
			o0 => And22580_o0
		);
		Nor22600 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i3,
			o0 => Nor22600_o0
		);
		And22620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22600_o0,
			i1 => Nor22060_o0,
			o0 => And22620_o0
		);
		And22640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22620_o0,
			i1 => And22580_o0,
			o0 => And22640_o0
		);
		And22660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22640_o0,
			i1 => Or22540_o0,
			o0 => And22660_o0
		);
		Or22680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22660_o0,
			i1 => And22200_o0,
			o0 => Or22680_o0
		);
		And22700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22680_o0,
			i1 => Not60_o0,
			o0 => And22700_o0
		);
		Nand22720 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i4,
			o0 => Nand22720_o0
		);
		And22740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand22720_o0,
			i1 => Not140_o0,
			o0 => And22740_o0
		);
		And22760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => i3,
			o0 => And22760_o0
		);
		Or22780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22760_o0,
			i1 => And22740_o0,
			o0 => Or22780_o0
		);
		And22800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i15,
			o0 => And22800_o0
		);
		And22820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22800_o0,
			i1 => Nor21220_o0,
			o0 => And22820_o0
		);
		Or22840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22820_o0,
			i1 => And22320_o0,
			o0 => Or22840_o0
		);
		And22860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22840_o0,
			i1 => i16,
			o0 => And22860_o0
		);
		And22880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22860_o0,
			i1 => Or22780_o0,
			o0 => And22880_o0
		);
		Nor22900 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i16,
			o0 => Nor22900_o0
		);
		And22920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22900_o0,
			i1 => And21100_o0,
			o0 => And22920_o0
		);
		And22940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not540_o0,
			o0 => And22940_o0
		);
		And22960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22940_o0,
			i1 => Nor22600_o0,
			o0 => And22960_o0
		);
		And22980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22960_o0,
			i1 => And22920_o0,
			o0 => And22980_o0
		);
		Or23000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22980_o0,
			i1 => And22880_o0,
			o0 => Or23000_o0
		);
		And23020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => Not180_o0,
			o0 => And23020_o0
		);
		And23040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Or23000_o0,
			o0 => And23040_o0
		);
		And23060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => And21820_o0,
			o0 => And23060_o0
		);
		And23080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not2080_o0,
			i1 => i12,
			o0 => And23080_o0
		);
		And23100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Not540_o0,
			o0 => And23100_o0
		);
		And23120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23100_o0,
			i1 => Nor22600_o0,
			o0 => And23120_o0
		);
		And23140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23120_o0,
			i1 => And23060_o0,
			o0 => And23140_o0
		);
		Or23160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23140_o0,
			i1 => And23040_o0,
			o0 => Or23160_o0
		);
		And23180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not100_o0,
			i1 => i0,
			o0 => And23180_o0
		);
		Nor23200 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i2,
			o0 => Nor23200_o0
		);
		And23220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23200_o0,
			i1 => And23180_o0,
			o0 => And23220_o0
		);
		And23240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23220_o0,
			i1 => Or23160_o0,
			o0 => And23240_o0
		);
		Or23260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23240_o0,
			i1 => And22700_o0,
			o0 => Or23260_o0
		);
		Nor23280 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i9,
			i1 => i8,
			o0 => Nor23280_o0
		);
		Not3300 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			o0 => Not3300_o0
		);
		Nor23320 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			i1 => i10,
			o0 => Nor23320_o0
		);
		And23340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23320_o0,
			i1 => Not3300_o0,
			o0 => And23340_o0
		);
		And23360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23340_o0,
			i1 => Nor23280_o0,
			o0 => And23360_o0
		);
		And23380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23360_o0,
			i1 => Or23260_o0,
			o0 => And23380_o0
		);
		And23400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22300_o0,
			i1 => And21100_o0,
			o0 => And23400_o0
		);
		Or23420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23400_o0,
			i1 => And22800_o0,
			o0 => Or23420_o0
		);
		And23440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1280_o0,
			i1 => i13,
			o0 => And23440_o0
		);
		And23460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23440_o0,
			i1 => Or23420_o0,
			o0 => And23460_o0
		);
		Or23480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23460_o0,
			i1 => Not2080_o0,
			o0 => Or23480_o0
		);
		And23500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or23480_o0,
			i1 => i14,
			o0 => And23500_o0
		);
		And23520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i13,
			o0 => And23520_o0
		);
		Nor23540 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i28,
			i1 => i15,
			o0 => Nor23540_o0
		);
		And23560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23540_o0,
			i1 => And23520_o0,
			o0 => And23560_o0
		);
		Or23580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23560_o0,
			i1 => And23500_o0,
			o0 => Or23580_o0
		);
		Nor23600 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i1,
			i1 => i0,
			o0 => Nor23600_o0
		);
		And23620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Nor21140_o0,
			o0 => And23620_o0
		);
		And23640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23620_o0,
			i1 => Nor23600_o0,
			o0 => And23640_o0
		);
		And23660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not3300_o0,
			i1 => i12,
			o0 => And23660_o0
		);
		And23680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23660_o0,
			i1 => i40,
			o0 => And23680_o0
		);
		And23700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23320_o0,
			i1 => Nor23280_o0,
			o0 => And23700_o0
		);
		And23720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23700_o0,
			i1 => And23680_o0,
			o0 => And23720_o0
		);
		And23740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23720_o0,
			i1 => And23640_o0,
			o0 => And23740_o0
		);
		And23760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23740_o0,
			i1 => Or23580_o0,
			o0 => And23760_o0
		);
		And23780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22900_o0,
			i1 => i15,
			o0 => And23780_o0
		);
		Or23800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23780_o0,
			i1 => Not2080_o0,
			o0 => Or23800_o0
		);
		And23820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or23800_o0,
			i1 => i14,
			o0 => And23820_o0
		);
		Not3840 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i28,
			o0 => Not3840_o0
		);
		Nand23860 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i25,
			i1 => i24,
			o0 => Nand23860_o0
		);
		Or23880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand23860_o0,
			i1 => Not3840_o0,
			o0 => Or23880_o0
		);
		And23900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => Not620_o0,
			o0 => And23900_o0
		);
		And23920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23900_o0,
			i1 => Or23880_o0,
			o0 => And23920_o0
		);
		Or23940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And23920_o0,
			i1 => And23820_o0,
			o0 => Or23940_o0
		);
		And23960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or23940_o0,
			i1 => And23740_o0,
			o0 => And23960_o0
		);
		Or23980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i3,
			i1 => i2,
			o0 => Or23980_o0
		);
		Nor24000 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i12,
			o0 => Nor24000_o0
		);
		And24020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24000_o0,
			i1 => Or23980_o0,
			o0 => And24020_o0
		);
		And24040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i14,
			o0 => And24040_o0
		);
		And24060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24040_o0,
			i1 => i12,
			o0 => And24060_o0
		);
		And24080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24060_o0,
			i1 => Nor21140_o0,
			o0 => And24080_o0
		);
		Or24100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24080_o0,
			i1 => And24020_o0,
			o0 => Or24100_o0
		);
		And24120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24100_o0,
			i1 => Not1080_o0,
			o0 => And24120_o0
		);
		And24140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => Not140_o0,
			o0 => And24140_o0
		);
		And24160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24140_o0,
			i1 => Not120_o0,
			o0 => And24160_o0
		);
		And24180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i18,
			o0 => And24180_o0
		);
		And24200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24180_o0,
			i1 => i14,
			o0 => And24200_o0
		);
		And24220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24200_o0,
			i1 => And24160_o0,
			o0 => And24220_o0
		);
		Or24240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24220_o0,
			i1 => And24120_o0,
			o0 => Or24240_o0
		);
		And24260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24240_o0,
			i1 => Not540_o0,
			o0 => And24260_o0
		);
		And24280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not180_o0,
			i1 => i5,
			o0 => And24280_o0
		);
		Nor24300 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i14,
			o0 => Nor24300_o0
		);
		And24320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24300_o0,
			i1 => And24280_o0,
			o0 => And24320_o0
		);
		And24340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24320_o0,
			i1 => Or23980_o0,
			o0 => And24340_o0
		);
		Or24360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24340_o0,
			i1 => And24260_o0,
			o0 => Or24360_o0
		);
		And24380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24360_o0,
			i1 => Not160_o0,
			o0 => And24380_o0
		);
		And24400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => Not140_o0,
			o0 => And24400_o0
		);
		And24420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24400_o0,
			i1 => Not120_o0,
			o0 => And24420_o0
		);
		Or24440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24420_o0,
			i1 => Or23980_o0,
			o0 => Or24440_o0
		);
		And24460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not180_o0,
			i1 => i4,
			o0 => And24460_o0
		);
		And24480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24460_o0,
			i1 => Nor24300_o0,
			o0 => And24480_o0
		);
		And24500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24480_o0,
			i1 => Or24440_o0,
			o0 => And24500_o0
		);
		Or24520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24500_o0,
			i1 => And24380_o0,
			o0 => Or24520_o0
		);
		And24540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24520_o0,
			i1 => Not1280_o0,
			o0 => And24540_o0
		);
		And24560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i4,
			o0 => And24560_o0
		);
		And24580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24560_o0,
			i1 => Nor21140_o0,
			o0 => And24580_o0
		);
		Or24600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24580_o0,
			i1 => Or23980_o0,
			o0 => Or24600_o0
		);
		And24620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1080_o0,
			i1 => i16,
			o0 => And24620_o0
		);
		And24640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24620_o0,
			i1 => Nor24000_o0,
			o0 => And24640_o0
		);
		And24660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24640_o0,
			i1 => Or24600_o0,
			o0 => And24660_o0
		);
		Or24680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24660_o0,
			i1 => And24540_o0,
			o0 => Or24680_o0
		);
		And24700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24680_o0,
			i1 => Not100_o0,
			o0 => And24700_o0
		);
		Or24720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not540_o0,
			o0 => Or24720_o0
		);
		And24740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23200_o0,
			i1 => Not1080_o0,
			o0 => And24740_o0
		);
		And24760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22600_o0,
			i1 => And21420_o0,
			o0 => And24760_o0
		);
		And24780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24760_o0,
			i1 => And24740_o0,
			o0 => And24780_o0
		);
		And24800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24780_o0,
			i1 => Or24720_o0,
			o0 => And24800_o0
		);
		Or24820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24800_o0,
			i1 => And24700_o0,
			o0 => Or24820_o0
		);
		And24840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24820_o0,
			i1 => i15,
			o0 => And24840_o0
		);
		And24860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not140_o0,
			o0 => And24860_o0
		);
		And24880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not180_o0,
			o0 => And24880_o0
		);
		And24900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24880_o0,
			i1 => Nor22060_o0,
			o0 => And24900_o0
		);
		Nor24920 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i14,
			o0 => Nor24920_o0
		);
		And24940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not1080_o0,
			o0 => And24940_o0
		);
		And24960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24940_o0,
			i1 => Nor24920_o0,
			o0 => And24960_o0
		);
		And24980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24960_o0,
			i1 => And24900_o0,
			o0 => And24980_o0
		);
		And25000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24980_o0,
			i1 => And24860_o0,
			o0 => And25000_o0
		);
		And25020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => Not140_o0,
			o0 => And25020_o0
		);
		And25040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25020_o0,
			i1 => Not120_o0,
			o0 => And25040_o0
		);
		Or25060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25040_o0,
			i1 => Or23980_o0,
			o0 => Or25060_o0
		);
		And25080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25060_o0,
			i1 => i1,
			o0 => And25080_o0
		);
		Nor25100 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i1,
			o0 => Nor25100_o0
		);
		And25120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor25100_o0,
			i1 => And2560_o0,
			o0 => And25120_o0
		);
		And25140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25120_o0,
			i1 => Nor21140_o0,
			o0 => And25140_o0
		);
		Or25160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25140_o0,
			i1 => And25080_o0,
			o0 => Or25160_o0
		);
		And25180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25160_o0,
			i1 => Xor2960_o0,
			o0 => And25180_o0
		);
		Xor25200 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i4,
			o0 => Xor25200_o0
		);
		Xor25220 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i16,
			o0 => Xor25220_o0
		);
		Nor25240 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor25220_o0,
			i1 => i1,
			o0 => Nor25240_o0
		);
		And25260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor25240_o0,
			i1 => Xor25200_o0,
			o0 => And25260_o0
		);
		And25280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not1280_o0,
			o0 => And25280_o0
		);
		And25300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not160_o0,
			i1 => i1,
			o0 => And25300_o0
		);
		And25320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25300_o0,
			i1 => i5,
			o0 => And25320_o0
		);
		And25340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25320_o0,
			i1 => And25280_o0,
			o0 => And25340_o0
		);
		Or25360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25340_o0,
			i1 => And25260_o0,
			o0 => Or25360_o0
		);
		And25380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25360_o0,
			i1 => Nor21140_o0,
			o0 => And25380_o0
		);
		Or25400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25380_o0,
			i1 => And25180_o0,
			o0 => Or25400_o0
		);
		And25420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1080_o0,
			i1 => i15,
			o0 => And25420_o0
		);
		And25440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25420_o0,
			i1 => Nor24000_o0,
			o0 => And25440_o0
		);
		And25460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25440_o0,
			i1 => Or25400_o0,
			o0 => And25460_o0
		);
		Or25480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25460_o0,
			i1 => And25000_o0,
			o0 => Or25480_o0
		);
		Or25500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or25480_o0,
			i1 => And24840_o0,
			o0 => Or25500_o0
		);
		And25520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25500_o0,
			i1 => Not1040_o0,
			o0 => And25520_o0
		);
		Or25540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i3,
			o0 => Or25540_o0
		);
		Or25560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or25540_o0,
			i1 => i2,
			o0 => Or25560_o0
		);
		And25580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25560_o0,
			i1 => And2640_o0,
			o0 => And25580_o0
		);
		And25600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not1280_o0,
			o0 => And25600_o0
		);
		And25620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21140_o0,
			i1 => i15,
			o0 => And25620_o0
		);
		And25640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25620_o0,
			i1 => And25600_o0,
			o0 => And25640_o0
		);
		Or25660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25640_o0,
			i1 => And25580_o0,
			o0 => Or25660_o0
		);
		And25680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not180_o0,
			o0 => And25680_o0
		);
		And25700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25680_o0,
			i1 => And2240_o0,
			o0 => And25700_o0
		);
		And25720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25700_o0,
			i1 => Or25660_o0,
			o0 => And25720_o0
		);
		And25740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => Not620_o0,
			o0 => And25740_o0
		);
		And25760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2400_o0,
			i1 => i27,
			o0 => And25760_o0
		);
		And25780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25760_o0,
			i1 => And25740_o0,
			o0 => And25780_o0
		);
		And25800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i29,
			i1 => i15,
			o0 => And25800_o0
		);
		Or25820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25800_o0,
			i1 => And25780_o0,
			o0 => Or25820_o0
		);
		And25840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i12,
			o0 => And25840_o0
		);
		And25860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25840_o0,
			i1 => Nor21140_o0,
			o0 => And25860_o0
		);
		And25880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25860_o0,
			i1 => Or25820_o0,
			o0 => And25880_o0
		);
		Or25900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25880_o0,
			i1 => And25720_o0,
			o0 => Or25900_o0
		);
		And25920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25900_o0,
			i1 => Not100_o0,
			o0 => And25920_o0
		);
		And25940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2260_o0,
			i1 => i16,
			o0 => And25940_o0
		);
		And25960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21420_o0,
			i1 => Not620_o0,
			o0 => And25960_o0
		);
		And25980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25960_o0,
			i1 => And25940_o0,
			o0 => And25980_o0
		);
		Or26000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25980_o0,
			i1 => And25920_o0,
			o0 => Or26000_o0
		);
		And26020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26000_o0,
			i1 => Not540_o0,
			o0 => And26020_o0
		);
		And26040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i3,
			i1 => Not120_o0,
			o0 => And26040_o0
		);
		And26060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26040_o0,
			i1 => Not100_o0,
			o0 => And26060_o0
		);
		Or26080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i2,
			i1 => i1,
			o0 => Or26080_o0
		);
		Or26100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or26080_o0,
			i1 => And26060_o0,
			o0 => Or26100_o0
		);
		And26120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => i19,
			o0 => And26120_o0
		);
		And26140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24280_o0,
			i1 => And2640_o0,
			o0 => And26140_o0
		);
		And26160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26140_o0,
			i1 => And26120_o0,
			o0 => And26160_o0
		);
		And26180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26160_o0,
			i1 => Or26100_o0,
			o0 => And26180_o0
		);
		Or26200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26180_o0,
			i1 => And26020_o0,
			o0 => Or26200_o0
		);
		And26220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26200_o0,
			i1 => Not160_o0,
			o0 => And26220_o0
		);
		And26240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24400_o0,
			i1 => Nor22060_o0,
			o0 => And26240_o0
		);
		Or26260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26240_o0,
			i1 => Or26100_o0,
			o0 => Or26260_o0
		);
		And26280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24460_o0,
			i1 => And2640_o0,
			o0 => And26280_o0
		);
		And26300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26280_o0,
			i1 => And26120_o0,
			o0 => And26300_o0
		);
		And26320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26300_o0,
			i1 => Or26260_o0,
			o0 => And26320_o0
		);
		Or26340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26320_o0,
			i1 => And26220_o0,
			o0 => Or26340_o0
		);
		And26360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26340_o0,
			i1 => Not80_o0,
			o0 => And26360_o0
		);
		Or26380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26360_o0,
			i1 => And25520_o0,
			o0 => Or26380_o0
		);
		And26400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26380_o0,
			i1 => Not60_o0,
			o0 => And26400_o0
		);
		And26420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23200_o0,
			i1 => Not180_o0,
			o0 => And26420_o0
		);
		And26440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26420_o0,
			i1 => And23180_o0,
			o0 => And26440_o0
		);
		And26460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26440_o0,
			i1 => Or23000_o0,
			o0 => And26460_o0
		);
		Or26480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26460_o0,
			i1 => And26400_o0,
			o0 => Or26480_o0
		);
		And26500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26480_o0,
			i1 => i13,
			o0 => And26500_o0
		);
		And26520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not140_o0,
			o0 => And26520_o0
		);
		Xor26540 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i16,
			o0 => Xor26540_o0
		);
		Nor26560 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor26540_o0,
			i1 => i15,
			o0 => Nor26560_o0
		);
		And26580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => Not1280_o0,
			o0 => And26580_o0
		);
		And26600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26580_o0,
			i1 => i15,
			o0 => And26600_o0
		);
		Or26620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26600_o0,
			i1 => Nor26560_o0,
			o0 => Or26620_o0
		);
		And26640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26620_o0,
			i1 => And26520_o0,
			o0 => And26640_o0
		);
		Nor26660 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i16,
			o0 => Nor26660_o0
		);
		And26680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not620_o0,
			i1 => i3,
			o0 => And26680_o0
		);
		And26700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26680_o0,
			i1 => Nor26660_o0,
			o0 => And26700_o0
		);
		Or26720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26700_o0,
			i1 => And26640_o0,
			o0 => Or26720_o0
		);
		And26740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26720_o0,
			i1 => Not60_o0,
			o0 => And26740_o0
		);
		And26760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not140_o0,
			i1 => i0,
			o0 => And26760_o0
		);
		And26780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor26660_o0,
			i1 => Not620_o0,
			o0 => And26780_o0
		);
		And26800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26780_o0,
			i1 => And26760_o0,
			o0 => And26800_o0
		);
		Or26820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26800_o0,
			i1 => And26740_o0,
			o0 => Or26820_o0
		);
		And26840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26820_o0,
			i1 => And21520_o0,
			o0 => And26840_o0
		);
		And26860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Not80_o0,
			o0 => And26860_o0
		);
		And26880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22060_o0,
			i1 => Nor21260_o0,
			o0 => And26880_o0
		);
		And26900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26880_o0,
			i1 => And26860_o0,
			o0 => And26900_o0
		);
		And26920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26900_o0,
			i1 => And26840_o0,
			o0 => And26920_o0
		);
		Or26940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26920_o0,
			i1 => And26500_o0,
			o0 => Or26940_o0
		);
		And26960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or26940_o0,
			i1 => And23360_o0,
			o0 => And26960_o0
		);
		Xor26980 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i17,
			o0 => Xor26980_o0
		);
		Not7000 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Xor26980_o0,
			o0 => Not7000_o0
		);
		And27020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor2200_o0,
			i1 => i19,
			o0 => And27020_o0
		);
		And27040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27020_o0,
			i1 => Not7000_o0,
			o0 => And27040_o0
		);
		And27060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21240_o0,
			i1 => i16,
			o0 => And27060_o0
		);
		Or27080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27060_o0,
			i1 => And27040_o0,
			o0 => Or27080_o0
		);
		And27100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27080_o0,
			i1 => Not180_o0,
			o0 => And27100_o0
		);
		Not7120 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			o0 => Not7120_o0
		);
		Not7140 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i25,
			o0 => Not7140_o0
		);
		Or27160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => Not7140_o0,
			o0 => Or27160_o0
		);
		Or27180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or27160_o0,
			i1 => Not7120_o0,
			o0 => Or27180_o0
		);
		Or27200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or27180_o0,
			i1 => Not3840_o0,
			o0 => Or27200_o0
		);
		And27220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27200_o0,
			i1 => Not620_o0,
			o0 => And27220_o0
		);
		Or27240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27220_o0,
			i1 => And25800_o0,
			o0 => Or27240_o0
		);
		And27260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27240_o0,
			i1 => i12,
			o0 => And27260_o0
		);
		Or27280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27260_o0,
			i1 => And27100_o0,
			o0 => Or27280_o0
		);
		And27300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27280_o0,
			i1 => And26520_o0,
			o0 => And27300_o0
		);
		Or27320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27300_o0,
			i1 => And2840_o0,
			o0 => Or27320_o0
		);
		And27340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27320_o0,
			i1 => Not120_o0,
			o0 => And27340_o0
		);
		Or27360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27340_o0,
			i1 => And2900_o0,
			o0 => Or27360_o0
		);
		And27380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27360_o0,
			i1 => Not540_o0,
			o0 => And27380_o0
		);
		And27400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21020_o0,
			i1 => i3,
			o0 => And27400_o0
		);
		And27420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27400_o0,
			i1 => Not120_o0,
			o0 => And27420_o0
		);
		Not7440 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Xor25220_o0,
			o0 => Not7440_o0
		);
		And27460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor2960_o0,
			i1 => i2,
			o0 => And27460_o0
		);
		Or27480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27460_o0,
			i1 => Not7440_o0,
			o0 => Or27480_o0
		);
		And27500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22800_o0,
			i1 => Not1080_o0,
			o0 => And27500_o0
		);
		And27520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27500_o0,
			i1 => Or27480_o0,
			o0 => And27520_o0
		);
		And27540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => i2,
			o0 => And27540_o0
		);
		And27560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27540_o0,
			i1 => And2260_o0,
			o0 => And27560_o0
		);
		Or27580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27560_o0,
			i1 => And27520_o0,
			o0 => Or27580_o0
		);
		Or27600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or27580_o0,
			i1 => And27420_o0,
			o0 => Or27600_o0
		);
		And27620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27600_o0,
			i1 => And24280_o0,
			o0 => And27620_o0
		);
		Or27640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27620_o0,
			i1 => And27380_o0,
			o0 => Or27640_o0
		);
		And27660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27640_o0,
			i1 => Not160_o0,
			o0 => And27660_o0
		);
		And27680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21140_o0,
			i1 => i5,
			o0 => And27680_o0
		);
		And27700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27680_o0,
			i1 => Or21020_o0,
			o0 => And27700_o0
		);
		Or27720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27700_o0,
			i1 => Or27600_o0,
			o0 => Or27720_o0
		);
		And27740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27720_o0,
			i1 => And24460_o0,
			o0 => And27740_o0
		);
		Or27760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27740_o0,
			i1 => And27660_o0,
			o0 => Or27760_o0
		);
		And27780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27760_o0,
			i1 => Not100_o0,
			o0 => And27780_o0
		);
		Or27800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27780_o0,
			i1 => And21440_o0,
			o0 => Or27800_o0
		);
		And27820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27800_o0,
			i1 => Not60_o0,
			o0 => And27820_o0
		);
		Nor27840 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i2,
			o0 => Nor27840_o0
		);
		And27860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor27840_o0,
			i1 => And23180_o0,
			o0 => And27860_o0
		);
		And27880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27860_o0,
			i1 => Or23000_o0,
			o0 => And27880_o0
		);
		Or27900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27880_o0,
			i1 => And27820_o0,
			o0 => Or27900_o0
		);
		And27920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or27900_o0,
			i1 => i13,
			o0 => And27920_o0
		);
		And27940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Nor21260_o0,
			o0 => And27940_o0
		);
		And27960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27940_o0,
			i1 => Nor22060_o0,
			o0 => And27960_o0
		);
		And27980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27960_o0,
			i1 => And26840_o0,
			o0 => And27980_o0
		);
		Or28000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And27980_o0,
			i1 => And27920_o0,
			o0 => Or28000_o0
		);
		And28020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28000_o0,
			i1 => Not80_o0,
			o0 => And28020_o0
		);
		And28040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not1040_o0,
			o0 => And28040_o0
		);
		And28060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i14,
			o0 => And28060_o0
		);
		And28080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28060_o0,
			i1 => Not1280_o0,
			o0 => And28080_o0
		);
		And28100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28080_o0,
			i1 => And28040_o0,
			o0 => And28100_o0
		);
		And28120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => i12,
			o0 => And28120_o0
		);
		And28140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => Nor21260_o0,
			o0 => And28140_o0
		);
		And28160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23600_o0,
			i1 => Nor21140_o0,
			o0 => And28160_o0
		);
		And28180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28160_o0,
			i1 => And28140_o0,
			o0 => And28180_o0
		);
		And28200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28180_o0,
			i1 => And28100_o0,
			o0 => And28200_o0
		);
		Or28220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28200_o0,
			i1 => And28020_o0,
			o0 => Or28220_o0
		);
		And28240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28220_o0,
			i1 => And23360_o0,
			o0 => And28240_o0
		);
		And28260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => And21300_o0,
			o0 => And28260_o0
		);
		And28280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => And2640_o0,
			o0 => And28280_o0
		);
		Or28300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28280_o0,
			i1 => And28260_o0,
			o0 => Or28300_o0
		);
		And28320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28300_o0,
			i1 => i40,
			o0 => And28320_o0
		);
		And28340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28320_o0,
			i1 => Not540_o0,
			o0 => And28340_o0
		);
		And28360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => And2640_o0,
			o0 => And28360_o0
		);
		Or28380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28360_o0,
			i1 => And2600_o0,
			o0 => Or28380_o0
		);
		And28400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28380_o0,
			i1 => i5,
			o0 => And28400_o0
		);
		Or28420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28400_o0,
			i1 => And28340_o0,
			o0 => Or28420_o0
		);
		And28440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28420_o0,
			i1 => i19,
			o0 => And28440_o0
		);
		And28460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i5,
			o0 => And28460_o0
		);
		And28480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i16,
			o0 => And28480_o0
		);
		And28500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28480_o0,
			i1 => Nor21980_o0,
			o0 => And28500_o0
		);
		Or28520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28500_o0,
			i1 => And28460_o0,
			o0 => Or28520_o0
		);
		And28540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => Not1500_o0,
			o0 => And28540_o0
		);
		And28560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28540_o0,
			i1 => Or28520_o0,
			o0 => And28560_o0
		);
		Or28580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28560_o0,
			i1 => And28440_o0,
			o0 => Or28580_o0
		);
		And28600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28580_o0,
			i1 => Not180_o0,
			o0 => And28600_o0
		);
		And28620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => i12,
			o0 => And28620_o0
		);
		And28640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28620_o0,
			i1 => Or27240_o0,
			o0 => And28640_o0
		);
		Or28660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28640_o0,
			i1 => And28600_o0,
			o0 => Or28660_o0
		);
		And28680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28660_o0,
			i1 => Not160_o0,
			o0 => And28680_o0
		);
		Or28700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28680_o0,
			i1 => And2780_o0,
			o0 => Or28700_o0
		);
		And28720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28700_o0,
			i1 => Not140_o0,
			o0 => And28720_o0
		);
		Or28740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28720_o0,
			i1 => And2840_o0,
			o0 => Or28740_o0
		);
		And28760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28740_o0,
			i1 => Not120_o0,
			o0 => And28760_o0
		);
		Or28780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28760_o0,
			i1 => And2900_o0,
			o0 => Or28780_o0
		);
		And28800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28780_o0,
			i1 => Not100_o0,
			o0 => And28800_o0
		);
		Or28820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28800_o0,
			i1 => And21440_o0,
			o0 => Or28820_o0
		);
		And28840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28820_o0,
			i1 => Not60_o0,
			o0 => And28840_o0
		);
		And28860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22840_o0,
			i1 => Nand22720_o0,
			o0 => And28860_o0
		);
		And28880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28860_o0,
			i1 => i16,
			o0 => And28880_o0
		);
		And28900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22940_o0,
			i1 => Not160_o0,
			o0 => And28900_o0
		);
		And28920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28900_o0,
			i1 => And22920_o0,
			o0 => And28920_o0
		);
		Or28940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28920_o0,
			i1 => And28880_o0,
			o0 => Or28940_o0
		);
		And28960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21140_o0,
			i1 => Not180_o0,
			o0 => And28960_o0
		);
		And28980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28960_o0,
			i1 => And23180_o0,
			o0 => And28980_o0
		);
		And29000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28980_o0,
			i1 => Or28940_o0,
			o0 => And29000_o0
		);
		Or29020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29000_o0,
			i1 => And28840_o0,
			o0 => Or29020_o0
		);
		And29040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29020_o0,
			i1 => Not80_o0,
			o0 => And29040_o0
		);
		And29060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => i12,
			o0 => And29060_o0
		);
		And29080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29060_o0,
			i1 => And28160_o0,
			o0 => And29080_o0
		);
		And29100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29080_o0,
			i1 => And28100_o0,
			o0 => And29100_o0
		);
		Or29120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29100_o0,
			i1 => And29040_o0,
			o0 => Or29120_o0
		);
		And29140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29120_o0,
			i1 => i13,
			o0 => And29140_o0
		);
		And29160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => i18,
			o0 => And29160_o0
		);
		And29180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29160_o0,
			i1 => Xor2200_o0,
			o0 => And29180_o0
		);
		And29200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not620_o0,
			i1 => i5,
			o0 => And29200_o0
		);
		And29220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29200_o0,
			i1 => Nor26660_o0,
			o0 => And29220_o0
		);
		Or29240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29220_o0,
			i1 => And29180_o0,
			o0 => Or29240_o0
		);
		Nor29260 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i13,
			o0 => Nor29260_o0
		);
		And29280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => And21520_o0,
			o0 => And29280_o0
		);
		And29300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22100_o0,
			i1 => Nor21140_o0,
			o0 => And29300_o0
		);
		And29320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29300_o0,
			i1 => Nor23600_o0,
			o0 => And29320_o0
		);
		And29340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29320_o0,
			i1 => And29280_o0,
			o0 => And29340_o0
		);
		And29360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29340_o0,
			i1 => Or29240_o0,
			o0 => And29360_o0
		);
		Or29380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29360_o0,
			i1 => And29140_o0,
			o0 => Or29380_o0
		);
		And29400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29380_o0,
			i1 => And23360_o0,
			o0 => And29400_o0
		);
		And29420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i32,
			i1 => i30,
			o0 => And29420_o0
		);
		And29440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29420_o0,
			i1 => i33,
			o0 => And29440_o0
		);
		Nor29460 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i31,
			i1 => i30,
			o0 => Nor29460_o0
		);
		Or29480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29460_o0,
			i1 => And29440_o0,
			o0 => Or29480_o0
		);
		And29500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29480_o0,
			i1 => i13,
			o0 => And29500_o0
		);
		And29520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => i17,
			o0 => And29520_o0
		);
		Not9540 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			o0 => Not9540_o0
		);
		And29560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			i1 => Not9540_o0,
			o0 => And29560_o0
		);
		Not9580 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			o0 => Not9580_o0
		);
		Or29600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not9580_o0,
			i1 => i26,
			o0 => Or29600_o0
		);
		And29620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29600_o0,
			i1 => i24,
			o0 => And29620_o0
		);
		Nor29640 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i24,
			o0 => Nor29640_o0
		);
		Or29660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29640_o0,
			i1 => And29620_o0,
			o0 => Or29660_o0
		);
		And29680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29660_o0,
			i1 => i23,
			o0 => And29680_o0
		);
		Not9700 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i23,
			o0 => Not9700_o0
		);
		And29720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9580_o0,
			i1 => i24,
			o0 => And29720_o0
		);
		And29740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29720_o0,
			i1 => Not9700_o0,
			o0 => And29740_o0
		);
		Or29760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29740_o0,
			i1 => And29680_o0,
			o0 => Or29760_o0
		);
		And29780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29760_o0,
			i1 => i22,
			o0 => And29780_o0
		);
		Not9800 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			o0 => Not9800_o0
		);
		And29820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29720_o0,
			i1 => Not9800_o0,
			o0 => And29820_o0
		);
		Or29840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29820_o0,
			i1 => And29780_o0,
			o0 => Or29840_o0
		);
		And29860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29840_o0,
			i1 => And29560_o0,
			o0 => And29860_o0
		);
		And29880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29860_o0,
			i1 => And29520_o0,
			o0 => And29880_o0
		);
		Or29900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29880_o0,
			i1 => Xor2200_o0,
			o0 => Or29900_o0
		);
		And29920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29900_o0,
			i1 => Not1500_o0,
			o0 => And29920_o0
		);
		And29940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not1040_o0,
			o0 => And29940_o0
		);
		And29960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29940_o0,
			i1 => And21300_o0,
			o0 => And29960_o0
		);
		Or29980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And29960_o0,
			i1 => And29920_o0,
			o0 => Or29980_o0
		);
		And210000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29980_o0,
			i1 => i18,
			o0 => And210000_o0
		);
		Nand210020 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i38,
			o0 => Nand210020_o0
		);
		And210040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210020_o0,
			i1 => Not1500_o0,
			o0 => And210040_o0
		);
		And210060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210040_o0,
			i1 => And2640_o0,
			o0 => And210060_o0
		);
		Or210080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210060_o0,
			i1 => And27020_o0,
			o0 => Or210080_o0
		);
		And210100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1080_o0,
			i1 => i17,
			o0 => And210100_o0
		);
		And210120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210100_o0,
			i1 => Or210080_o0,
			o0 => And210120_o0
		);
		Or210140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210120_o0,
			i1 => And210000_o0,
			o0 => Or210140_o0
		);
		And210160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210140_o0,
			i1 => Not2080_o0,
			o0 => And210160_o0
		);
		Or210180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210160_o0,
			i1 => And29500_o0,
			o0 => Or210180_o0
		);
		And210200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210180_o0,
			i1 => i12,
			o0 => And210200_o0
		);
		Xor210220 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i17,
			o0 => Xor210220_o0
		);
		And210240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => i19,
			o0 => And210240_o0
		);
		And210260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210240_o0,
			i1 => Xor210220_o0,
			o0 => And210260_o0
		);
		And210280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => i15,
			o0 => And210280_o0
		);
		Or210300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210280_o0,
			i1 => And28280_o0,
			o0 => Or210300_o0
		);
		Or210320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or210300_o0,
			i1 => And210260_o0,
			o0 => Or210320_o0
		);
		And210340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210320_o0,
			i1 => And23020_o0,
			o0 => And210340_o0
		);
		Or210360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210340_o0,
			i1 => And210200_o0,
			o0 => Or210360_o0
		);
		And210380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210360_o0,
			i1 => And2560_o0,
			o0 => And210380_o0
		);
		Or210400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i5,
			o0 => Or210400_o0
		);
		And210420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i16,
			o0 => And210420_o0
		);
		And210440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210420_o0,
			i1 => Not620_o0,
			o0 => And210440_o0
		);
		Or210460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210440_o0,
			i1 => And22800_o0,
			o0 => Or210460_o0
		);
		And210480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Not1080_o0,
			o0 => And210480_o0
		);
		And210500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210480_o0,
			i1 => Or210460_o0,
			o0 => And210500_o0
		);
		Not10520 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			o0 => Not10520_o0
		);
		And210540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not10520_o0,
			i1 => i20,
			o0 => And210540_o0
		);
		Nand210560 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i23,
			i1 => i22,
			o0 => Nand210560_o0
		);
		And210580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29560_o0,
			i1 => Not7120_o0,
			o0 => And210580_o0
		);
		And210600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210580_o0,
			i1 => Nand210560_o0,
			o0 => And210600_o0
		);
		Or210620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210600_o0,
			i1 => And210540_o0,
			o0 => Or210620_o0
		);
		Nand210640 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i26,
			i1 => i24,
			o0 => Nand210640_o0
		);
		And210660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210640_o0,
			i1 => i23,
			o0 => And210660_o0
		);
		And210680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => Not9700_o0,
			o0 => And210680_o0
		);
		Or210700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210680_o0,
			i1 => And210660_o0,
			o0 => Or210700_o0
		);
		And210720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210700_o0,
			i1 => i22,
			o0 => And210720_o0
		);
		And210740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => Not9800_o0,
			o0 => And210740_o0
		);
		Or210760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210740_o0,
			i1 => And210720_o0,
			o0 => Or210760_o0
		);
		And210780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29560_o0,
			i1 => i27,
			o0 => And210780_o0
		);
		And210800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210780_o0,
			i1 => Or210760_o0,
			o0 => And210800_o0
		);
		Or210820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210800_o0,
			i1 => Or210620_o0,
			o0 => Or210820_o0
		);
		And210840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210820_o0,
			i1 => i18,
			o0 => And210840_o0
		);
		And210860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29520_o0,
			i1 => And23080_o0,
			o0 => And210860_o0
		);
		And210880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210860_o0,
			i1 => And210840_o0,
			o0 => And210880_o0
		);
		Or210900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210880_o0,
			i1 => And210500_o0,
			o0 => Or210900_o0
		);
		And210920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210900_o0,
			i1 => Not1500_o0,
			o0 => And210920_o0
		);
		And210940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28380_o0,
			i1 => i19,
			o0 => And210940_o0
		);
		And210960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210940_o0,
			i1 => And23020_o0,
			o0 => And210960_o0
		);
		Or210980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210960_o0,
			i1 => And210920_o0,
			o0 => Or210980_o0
		);
		And211000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210980_o0,
			i1 => Or210400_o0,
			o0 => And211000_o0
		);
		And211020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i5,
			o0 => And211020_o0
		);
		Nor211040 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i13,
			o0 => Nor211040_o0
		);
		And211060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => And211020_o0,
			o0 => And211060_o0
		);
		And211080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211060_o0,
			i1 => And21960_o0,
			o0 => And211080_o0
		);
		Or211100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211080_o0,
			i1 => And211000_o0,
			o0 => Or211100_o0
		);
		Or211120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or211100_o0,
			i1 => And210380_o0,
			o0 => Or211120_o0
		);
		And211140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211120_o0,
			i1 => Not160_o0,
			o0 => And211140_o0
		);
		And211160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And2600_o0,
			o0 => And211160_o0
		);
		And211180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => Not1500_o0,
			o0 => And211180_o0
		);
		And211200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211180_o0,
			i1 => Or210620_o0,
			o0 => And211200_o0
		);
		And211220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211200_o0,
			i1 => And21640_o0,
			o0 => And211220_o0
		);
		And211240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Not620_o0,
			o0 => And211240_o0
		);
		And211260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211240_o0,
			i1 => And211220_o0,
			o0 => And211260_o0
		);
		Or211280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211260_o0,
			i1 => And211160_o0,
			o0 => Or211280_o0
		);
		And211300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211280_o0,
			i1 => Not1280_o0,
			o0 => And211300_o0
		);
		Or211320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And22320_o0,
			i1 => And2600_o0,
			o0 => Or211320_o0
		);
		And211340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => i16,
			o0 => And211340_o0
		);
		And211360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211340_o0,
			i1 => Or211320_o0,
			o0 => And211360_o0
		);
		Or211380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211360_o0,
			i1 => And211300_o0,
			o0 => Or211380_o0
		);
		And211400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211380_o0,
			i1 => i4,
			o0 => And211400_o0
		);
		Or211420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211400_o0,
			i1 => And211140_o0,
			o0 => Or211420_o0
		);
		And211440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211420_o0,
			i1 => Not140_o0,
			o0 => And211440_o0
		);
		And211460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Or2680_o0,
			o0 => And211460_o0
		);
		And211480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211460_o0,
			i1 => i3,
			o0 => And211480_o0
		);
		Or211500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211480_o0,
			i1 => And211440_o0,
			o0 => Or211500_o0
		);
		And211520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211500_o0,
			i1 => Not120_o0,
			o0 => And211520_o0
		);
		And211540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211460_o0,
			i1 => i2,
			o0 => And211540_o0
		);
		Or211560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211540_o0,
			i1 => And211520_o0,
			o0 => Or211560_o0
		);
		And211580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211560_o0,
			i1 => Not100_o0,
			o0 => And211580_o0
		);
		And211600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21420_o0,
			i1 => i13,
			o0 => And211600_o0
		);
		And211620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211600_o0,
			i1 => Or21400_o0,
			o0 => And211620_o0
		);
		Or211640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211620_o0,
			i1 => And211580_o0,
			o0 => Or211640_o0
		);
		And211660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211640_o0,
			i1 => Not60_o0,
			o0 => And211660_o0
		);
		And211680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28940_o0,
			i1 => And23020_o0,
			o0 => And211680_o0
		);
		And211700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27940_o0,
			i1 => And23060_o0,
			o0 => And211700_o0
		);
		Or211720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211700_o0,
			i1 => And211680_o0,
			o0 => Or211720_o0
		);
		And211740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23180_o0,
			i1 => Nor21140_o0,
			o0 => And211740_o0
		);
		And211760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211740_o0,
			i1 => Or211720_o0,
			o0 => And211760_o0
		);
		Or211780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211760_o0,
			i1 => And211660_o0,
			o0 => Or211780_o0
		);
		And211800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211780_o0,
			i1 => Not80_o0,
			o0 => And211800_o0
		);
		And211820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => And2640_o0,
			o0 => And211820_o0
		);
		Or211840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211820_o0,
			i1 => And26600_o0,
			o0 => Or211840_o0
		);
		And211860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i12,
			o0 => And211860_o0
		);
		And211880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211860_o0,
			i1 => Or211840_o0,
			o0 => And211880_o0
		);
		Or211900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211880_o0,
			i1 => Not180_o0,
			o0 => Or211900_o0
		);
		And211920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211900_o0,
			i1 => i13,
			o0 => And211920_o0
		);
		And211940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not2080_o0,
			o0 => And211940_o0
		);
		And211960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211940_o0,
			i1 => i12,
			o0 => And211960_o0
		);
		Or211980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And211960_o0,
			i1 => And211920_o0,
			o0 => Or211980_o0
		);
		And212000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24040_o0,
			i1 => Nor21260_o0,
			o0 => And212000_o0
		);
		And212020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212000_o0,
			i1 => And28160_o0,
			o0 => And212020_o0
		);
		And212040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212020_o0,
			i1 => Or211980_o0,
			o0 => And212040_o0
		);
		Or212060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212040_o0,
			i1 => And211800_o0,
			o0 => Or212060_o0
		);
		And212080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212060_o0,
			i1 => And23360_o0,
			o0 => And212080_o0
		);
		Not12100 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i8,
			o0 => Not12100_o0
		);
		Not12120 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			o0 => Not12120_o0
		);
		Or212140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			i1 => Not12120_o0,
			o0 => Or212140_o0
		);
		And212160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212140_o0,
			i1 => i9,
			o0 => And212160_o0
		);
		And212180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i16,
			o0 => And212180_o0
		);
		And212200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212180_o0,
			i1 => Not620_o0,
			o0 => And212200_o0
		);
		And212220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor26660_o0,
			i1 => i15,
			o0 => And212220_o0
		);
		Not12240 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i37,
			o0 => Not12240_o0
		);
		Nor212260 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i38,
			o0 => Nor212260_o0
		);
		And212280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => Not12240_o0,
			o0 => And212280_o0
		);
		And212300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212280_o0,
			i1 => And212220_o0,
			o0 => And212300_o0
		);
		Or212320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212300_o0,
			i1 => And212200_o0,
			o0 => Or212320_o0
		);
		And212340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212320_o0,
			i1 => And23080_o0,
			o0 => And212340_o0
		);
		And212360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And21300_o0,
			o0 => And212360_o0
		);
		And212380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12240_o0,
			i1 => i18,
			o0 => And212380_o0
		);
		And212400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212380_o0,
			i1 => Nor212260_o0,
			o0 => And212400_o0
		);
		And212420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212400_o0,
			i1 => And212360_o0,
			o0 => And212420_o0
		);
		Or212440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212420_o0,
			i1 => And212340_o0,
			o0 => Or212440_o0
		);
		And212460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212440_o0,
			i1 => Not1500_o0,
			o0 => And212460_o0
		);
		And212480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212280_o0,
			i1 => And2240_o0,
			o0 => And212480_o0
		);
		And212500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212480_o0,
			i1 => And212360_o0,
			o0 => And212500_o0
		);
		Or212520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212500_o0,
			i1 => And212460_o0,
			o0 => Or212520_o0
		);
		And212540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212520_o0,
			i1 => Not1040_o0,
			o0 => And212540_o0
		);
		And212560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210040_o0,
			i1 => Not1080_o0,
			o0 => And212560_o0
		);
		And212580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => And21740_o0,
			o0 => And212580_o0
		);
		And212600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212580_o0,
			i1 => And212560_o0,
			o0 => And212600_o0
		);
		Or212620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212600_o0,
			i1 => And212540_o0,
			o0 => Or212620_o0
		);
		Nor212640 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i11,
			o0 => Nor212640_o0
		);
		And212660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not3300_o0,
			o0 => And212660_o0
		);
		And212680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212660_o0,
			i1 => Nor212640_o0,
			o0 => And212680_o0
		);
		Nor212700 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => i9,
			o0 => Nor212700_o0
		);
		And212720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212700_o0,
			i1 => Nor21260_o0,
			o0 => And212720_o0
		);
		And212740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212720_o0,
			i1 => And28160_o0,
			o0 => And212740_o0
		);
		And212760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212740_o0,
			i1 => And212680_o0,
			o0 => And212760_o0
		);
		And212780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212760_o0,
			i1 => Or212620_o0,
			o0 => And212780_o0
		);
		Or212800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212780_o0,
			i1 => And212160_o0,
			o0 => Or212800_o0
		);
		And212820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212800_o0,
			i1 => Not12100_o0,
			o0 => And212820_o0
		);
		Not12840 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i30,
			o0 => Not12840_o0
		);
		And212860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => Not12840_o0,
			o0 => And212860_o0
		);
		And212880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => Not1040_o0,
			o0 => And212880_o0
		);
		And212900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => Not1280_o0,
			o0 => And212900_o0
		);
		And212920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212900_o0,
			i1 => i14,
			o0 => And212920_o0
		);
		Nor212940 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i30,
			i1 => i14,
			o0 => Nor212940_o0
		);
		Or212960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212940_o0,
			i1 => And212920_o0,
			o0 => Or212960_o0
		);
		And212980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or212960_o0,
			i1 => i15,
			o0 => And212980_o0
		);
		Or213000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212980_o0,
			i1 => And212860_o0,
			o0 => Or213000_o0
		);
		And213020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213000_o0,
			i1 => i13,
			o0 => And213020_o0
		);
		And213040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210100_o0,
			i1 => Nand210020_o0,
			o0 => And213040_o0
		);
		Or213060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213040_o0,
			i1 => And212880_o0,
			o0 => Or213060_o0
		);
		And213080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => Not1500_o0,
			o0 => And213080_o0
		);
		And213100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213080_o0,
			i1 => Nor29260_o0,
			o0 => And213100_o0
		);
		And213120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213100_o0,
			i1 => Or213060_o0,
			o0 => And213120_o0
		);
		Or213140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213120_o0,
			i1 => And213020_o0,
			o0 => Or213140_o0
		);
		And213160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213140_o0,
			i1 => i12,
			o0 => And213160_o0
		);
		And213180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not620_o0,
			i1 => i14,
			o0 => And213180_o0
		);
		And213200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => And23020_o0,
			o0 => And213200_o0
		);
		Or213220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213200_o0,
			i1 => And213160_o0,
			o0 => Or213220_o0
		);
		And213240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212660_o0,
			i1 => Nor23320_o0,
			o0 => And213240_o0
		);
		And213260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23280_o0,
			i1 => Nor21260_o0,
			o0 => And213260_o0
		);
		And213280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213260_o0,
			i1 => And28160_o0,
			o0 => And213280_o0
		);
		And213300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213280_o0,
			i1 => And213240_o0,
			o0 => And213300_o0
		);
		And213320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213300_o0,
			i1 => Or213220_o0,
			o0 => And213320_o0
		);
		Or213340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not1280_o0,
			i1 => i14,
			o0 => Or213340_o0
		);
		And213360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213340_o0,
			i1 => Not180_o0,
			o0 => And213360_o0
		);
		Nand213380 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i33,
			i1 => i32,
			o0 => Nand213380_o0
		);
		Or213400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand213380_o0,
			i1 => Not12840_o0,
			o0 => Or213400_o0
		);
		And213420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213400_o0,
			i1 => Not80_o0,
			o0 => And213420_o0
		);
		And213440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213420_o0,
			i1 => i12,
			o0 => And213440_o0
		);
		Or213460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213440_o0,
			i1 => And213360_o0,
			o0 => Or213460_o0
		);
		And213480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213460_o0,
			i1 => Not620_o0,
			o0 => And213480_o0
		);
		Or213500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213420_o0,
			i1 => And212920_o0,
			o0 => Or213500_o0
		);
		And213520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i12,
			o0 => And213520_o0
		);
		And213540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213520_o0,
			i1 => Or213500_o0,
			o0 => And213540_o0
		);
		Or213560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213540_o0,
			i1 => And213480_o0,
			o0 => Or213560_o0
		);
		And213580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213560_o0,
			i1 => i13,
			o0 => And213580_o0
		);
		And213600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213120_o0,
			i1 => i12,
			o0 => And213600_o0
		);
		Or213620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213600_o0,
			i1 => And213580_o0,
			o0 => Or213620_o0
		);
		And213640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213620_o0,
			i1 => And213300_o0,
			o0 => And213640_o0
		);
		Or213660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212400_o0,
			i1 => Not1080_o0,
			o0 => Or213660_o0
		);
		And213680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213660_o0,
			i1 => Nor24000_o0,
			o0 => And213680_o0
		);
		And213700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i14,
			o0 => And213700_o0
		);
		And213720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213700_o0,
			i1 => i12,
			o0 => And213720_o0
		);
		Or213740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213720_o0,
			i1 => And213680_o0,
			o0 => Or213740_o0
		);
		And213760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213740_o0,
			i1 => Not1280_o0,
			o0 => And213760_o0
		);
		Or213780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213760_o0,
			i1 => And24640_o0,
			o0 => Or213780_o0
		);
		And213800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213780_o0,
			i1 => Not1040_o0,
			o0 => And213800_o0
		);
		Not13820 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i33,
			o0 => Not13820_o0
		);
		Nor213840 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i35,
			i1 => Not13820_o0,
			o0 => Nor213840_o0
		);
		Nand213860 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => Nor213840_o0,
			i1 => i32,
			o0 => Nand213860_o0
		);
		Or213880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand213860_o0,
			i1 => Not12840_o0,
			o0 => Or213880_o0
		);
		And213900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i12,
			o0 => And213900_o0
		);
		And213920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213900_o0,
			i1 => Or213880_o0,
			o0 => And213920_o0
		);
		Or213940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And213920_o0,
			i1 => And213800_o0,
			o0 => Or213940_o0
		);
		And213960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213940_o0,
			i1 => i15,
			o0 => And213960_o0
		);
		And213980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213880_o0,
			i1 => i12,
			o0 => And213980_o0
		);
		And214000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24880_o0,
			i1 => And2260_o0,
			o0 => And214000_o0
		);
		Or214020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214000_o0,
			i1 => And213980_o0,
			o0 => Or214020_o0
		);
		And214040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214020_o0,
			i1 => Nor24920_o0,
			o0 => And214040_o0
		);
		Or214060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214040_o0,
			i1 => And213960_o0,
			o0 => Or214060_o0
		);
		And214080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214060_o0,
			i1 => i13,
			o0 => And214080_o0
		);
		And214100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i17,
			o0 => And214100_o0
		);
		Nor214120 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i17,
			o0 => Nor214120_o0
		);
		And214140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214120_o0,
			i1 => And212280_o0,
			o0 => And214140_o0
		);
		Or214160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214140_o0,
			i1 => And214100_o0,
			o0 => Or214160_o0
		);
		And214180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214160_o0,
			i1 => And21300_o0,
			o0 => And214180_o0
		);
		And214200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214100_o0,
			i1 => And2640_o0,
			o0 => And214200_o0
		);
		Or214220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214200_o0,
			i1 => And214180_o0,
			o0 => Or214220_o0
		);
		And214240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24300_o0,
			i1 => And23080_o0,
			o0 => And214240_o0
		);
		And214260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214240_o0,
			i1 => Or214220_o0,
			o0 => And214260_o0
		);
		Or214280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214260_o0,
			i1 => And214080_o0,
			o0 => Or214280_o0
		);
		And214300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214280_o0,
			i1 => And2560_o0,
			o0 => And214300_o0
		);
		And214320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Not1280_o0,
			o0 => And214320_o0
		);
		And214340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214320_o0,
			i1 => And210840_o0,
			o0 => And214340_o0
		);
		And214360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24620_o0,
			i1 => And23020_o0,
			o0 => And214360_o0
		);
		Or214380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214360_o0,
			i1 => And214340_o0,
			o0 => Or214380_o0
		);
		And214400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not80_o0,
			o0 => And214400_o0
		);
		And214420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214400_o0,
			i1 => Not1500_o0,
			o0 => And214420_o0
		);
		And214440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214420_o0,
			i1 => And29200_o0,
			o0 => And214440_o0
		);
		And214460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214440_o0,
			i1 => Or214380_o0,
			o0 => And214460_o0
		);
		Or214480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214460_o0,
			i1 => And214300_o0,
			o0 => Or214480_o0
		);
		And214500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214480_o0,
			i1 => Not160_o0,
			o0 => And214500_o0
		);
		And214520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211220_o0,
			i1 => Nor21840_o0,
			o0 => And214520_o0
		);
		And214540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214520_o0,
			i1 => And26860_o0,
			o0 => And214540_o0
		);
		And214560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214540_o0,
			i1 => i4,
			o0 => And214560_o0
		);
		Or214580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214560_o0,
			i1 => And214500_o0,
			o0 => Or214580_o0
		);
		And214600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214580_o0,
			i1 => Not60_o0,
			o0 => And214600_o0
		);
		And214620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not160_o0,
			i1 => i0,
			o0 => And214620_o0
		);
		And214640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214620_o0,
			i1 => And23100_o0,
			o0 => And214640_o0
		);
		And214660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => Not80_o0,
			o0 => And214660_o0
		);
		And214680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214660_o0,
			i1 => And21820_o0,
			o0 => And214680_o0
		);
		And214700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214680_o0,
			i1 => And214640_o0,
			o0 => And214700_o0
		);
		Or214720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214700_o0,
			i1 => And214600_o0,
			o0 => Or214720_o0
		);
		Nor214740 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i9,
			i1 => i3,
			o0 => Nor214740_o0
		);
		And214760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214740_o0,
			i1 => Nor22060_o0,
			o0 => And214760_o0
		);
		And214780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214760_o0,
			i1 => And23340_o0,
			o0 => And214780_o0
		);
		And214800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214780_o0,
			i1 => Or214720_o0,
			o0 => And214800_o0
		);
		Or214820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214800_o0,
			i1 => And212160_o0,
			o0 => Or214820_o0
		);
		And214840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214820_o0,
			i1 => Not12100_o0,
			o0 => And214840_o0
		);
		And214860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not540_o0,
			i1 => i4,
			o0 => And214860_o0
		);
		And214880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214540_o0,
			i1 => And214860_o0,
			o0 => And214880_o0
		);
		Or214900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214880_o0,
			i1 => And214500_o0,
			o0 => Or214900_o0
		);
		And214920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or214900_o0,
			i1 => Not60_o0,
			o0 => And214920_o0
		);
		Or214940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And214920_o0,
			i1 => And214700_o0,
			o0 => Or214940_o0
		);
		Nor214960 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => i8,
			o0 => Nor214960_o0
		);
		Nor214980 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i11,
			o0 => Nor214980_o0
		);
		And215000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214980_o0,
			i1 => Nor214960_o0,
			o0 => And215000_o0
		);
		And215020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215000_o0,
			i1 => And214760_o0,
			o0 => And215020_o0
		);
		And215040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215020_o0,
			i1 => Or214940_o0,
			o0 => And215040_o0
		);
		And215060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1500_o0,
			i1 => i18,
			o0 => And215060_o0
		);
		And215080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => Not1040_o0,
			o0 => And215080_o0
		);
		And215100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215080_o0,
			i1 => And2640_o0,
			o0 => And215100_o0
		);
		Or215120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215100_o0,
			i1 => And210120_o0,
			o0 => Or215120_o0
		);
		And215140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215120_o0,
			i1 => Not2080_o0,
			o0 => And215140_o0
		);
		And215160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or213880_o0,
			i1 => i13,
			o0 => And215160_o0
		);
		Or215180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215160_o0,
			i1 => And215140_o0,
			o0 => Or215180_o0
		);
		And215200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215180_o0,
			i1 => And2560_o0,
			o0 => And215200_o0
		);
		And215220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210820_o0,
			i1 => Not1500_o0,
			o0 => And215220_o0
		);
		And215240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215220_o0,
			i1 => And21640_o0,
			o0 => And215240_o0
		);
		Nor215260 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i13,
			o0 => Nor215260_o0
		);
		And215280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215260_o0,
			i1 => And29200_o0,
			o0 => And215280_o0
		);
		And215300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215280_o0,
			i1 => And215240_o0,
			o0 => And215300_o0
		);
		Or215320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215300_o0,
			i1 => And215200_o0,
			o0 => Or215320_o0
		);
		And215340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215320_o0,
			i1 => i12,
			o0 => And215340_o0
		);
		And215360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or211320_o0,
			i1 => And2560_o0,
			o0 => And215360_o0
		);
		And215380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29200_o0,
			i1 => And21820_o0,
			o0 => And215380_o0
		);
		Or215400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215380_o0,
			i1 => And215360_o0,
			o0 => Or215400_o0
		);
		And215420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215400_o0,
			i1 => i16,
			o0 => And215420_o0
		);
		And215440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24940_o0,
			i1 => Not1040_o0,
			o0 => And215440_o0
		);
		And215460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22940_o0,
			i1 => Not1280_o0,
			o0 => And215460_o0
		);
		And215480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215460_o0,
			i1 => And215440_o0,
			o0 => And215480_o0
		);
		Or215500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215480_o0,
			i1 => And215420_o0,
			o0 => Or215500_o0
		);
		And215520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215500_o0,
			i1 => And23020_o0,
			o0 => And215520_o0
		);
		Or215540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215520_o0,
			i1 => And215340_o0,
			o0 => Or215540_o0
		);
		And215560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215540_o0,
			i1 => Not160_o0,
			o0 => And215560_o0
		);
		And215580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24560_o0,
			i1 => And23080_o0,
			o0 => And215580_o0
		);
		And215600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215580_o0,
			i1 => And214520_o0,
			o0 => And215600_o0
		);
		Or215620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215600_o0,
			i1 => And215560_o0,
			o0 => Or215620_o0
		);
		And215640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215620_o0,
			i1 => Not60_o0,
			o0 => And215640_o0
		);
		And215660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214640_o0,
			i1 => And23060_o0,
			o0 => And215660_o0
		);
		Or215680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215660_o0,
			i1 => And215640_o0,
			o0 => Or215680_o0
		);
		Nor215700 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i14,
			o0 => Nor215700_o0
		);
		And215720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215700_o0,
			i1 => Nor23320_o0,
			o0 => And215720_o0
		);
		And215740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215720_o0,
			i1 => And214760_o0,
			o0 => And215740_o0
		);
		And215760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215740_o0,
			i1 => Or215680_o0,
			o0 => And215760_o0
		);
		Or215780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215760_o0,
			i1 => And212160_o0,
			o0 => Or215780_o0
		);
		And215800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215780_o0,
			i1 => Not12100_o0,
			o0 => And215800_o0
		);
		And215820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i16,
			o0 => And215820_o0
		);
		And215840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215820_o0,
			i1 => And214860_o0,
			o0 => And215840_o0
		);
		And215860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => Not160_o0,
			o0 => And215860_o0
		);
		Nor215880 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i16,
			o0 => Nor215880_o0
		);
		And215900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215880_o0,
			i1 => And215860_o0,
			o0 => And215900_o0
		);
		Or215920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215900_o0,
			i1 => And215840_o0,
			o0 => Or215920_o0
		);
		And215940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i1,
			o0 => And215940_o0
		);
		And215960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215940_o0,
			i1 => Or215920_o0,
			o0 => And215960_o0
		);
		And215980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28500_o0,
			i1 => Nor25100_o0,
			o0 => And215980_o0
		);
		Or216000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And215980_o0,
			i1 => And215960_o0,
			o0 => Or216000_o0
		);
		And216020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216000_o0,
			i1 => Not1080_o0,
			o0 => And216020_o0
		);
		And216040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24180_o0,
			i1 => i16,
			o0 => And216040_o0
		);
		And216060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216040_o0,
			i1 => Nor21980_o0,
			o0 => And216060_o0
		);
		And216080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216060_o0,
			i1 => Nor25100_o0,
			o0 => And216080_o0
		);
		Or216100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216080_o0,
			i1 => And216020_o0,
			o0 => Or216100_o0
		);
		And216120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216100_o0,
			i1 => Not1040_o0,
			o0 => And216120_o0
		);
		Xor216140 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i18,
			o0 => Xor216140_o0
		);
		And216160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor216140_o0,
			i1 => i17,
			o0 => And216160_o0
		);
		Or216180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216160_o0,
			i1 => Not1280_o0,
			o0 => Or216180_o0
		);
		And216200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216180_o0,
			i1 => Not620_o0,
			o0 => And216200_o0
		);
		And216220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2260_o0,
			i1 => And21300_o0,
			o0 => And216220_o0
		);
		Or216240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216220_o0,
			i1 => And216200_o0,
			o0 => Or216240_o0
		);
		And216260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216240_o0,
			i1 => And2560_o0,
			o0 => And216260_o0
		);
		And216280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => i5,
			o0 => And216280_o0
		);
		And216300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216280_o0,
			i1 => And21820_o0,
			o0 => And216300_o0
		);
		Or216320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216300_o0,
			i1 => And216260_o0,
			o0 => Or216320_o0
		);
		And216340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216320_o0,
			i1 => Nor25100_o0,
			o0 => And216340_o0
		);
		Or216360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216340_o0,
			i1 => And216120_o0,
			o0 => Or216360_o0
		);
		And216380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216360_o0,
			i1 => Not180_o0,
			o0 => And216380_o0
		);
		Nand216400 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i15,
			o0 => Nand216400_o0
		);
		And216420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28620_o0,
			i1 => Nor25100_o0,
			o0 => And216420_o0
		);
		And216440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216420_o0,
			i1 => Nand216400_o0,
			o0 => And216440_o0
		);
		Or216460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216440_o0,
			i1 => And216380_o0,
			o0 => Or216460_o0
		);
		And216480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216460_o0,
			i1 => i13,
			o0 => And216480_o0
		);
		And216500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i4,
			o0 => And216500_o0
		);
		And216520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216500_o0,
			i1 => And29940_o0,
			o0 => And216520_o0
		);
		And216540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			i1 => i20,
			o0 => And216540_o0
		);
		And216560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216540_o0,
			i1 => Not1500_o0,
			o0 => And216560_o0
		);
		And216580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22300_o0,
			i1 => Not160_o0,
			o0 => And216580_o0
		);
		And216600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216580_o0,
			i1 => And216560_o0,
			o0 => And216600_o0
		);
		Or216620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216600_o0,
			i1 => And216520_o0,
			o0 => Or216620_o0
		);
		And216640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216620_o0,
			i1 => i5,
			o0 => And216640_o0
		);
		And216660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214120_o0,
			i1 => Not620_o0,
			o0 => And216660_o0
		);
		Or216680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216660_o0,
			i1 => Xor21620_o0,
			o0 => Or216680_o0
		);
		And216700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => i40,
			o0 => And216700_o0
		);
		And216720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216700_o0,
			i1 => Or216680_o0,
			o0 => And216720_o0
		);
		Or216740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216720_o0,
			i1 => And216640_o0,
			o0 => Or216740_o0
		);
		And216760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216740_o0,
			i1 => i18,
			o0 => And216760_o0
		);
		Xor216780 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not620_o0,
			o0 => Xor216780_o0
		);
		Not16800 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i38,
			o0 => Not16800_o0
		);
		And216820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not16800_o0,
			i1 => i37,
			o0 => And216820_o0
		);
		Nand216840 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => And216820_o0,
			i1 => i39,
			o0 => Nand216840_o0
		);
		And216860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand216840_o0,
			i1 => And22300_o0,
			o0 => And216860_o0
		);
		Or216880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216860_o0,
			i1 => And22800_o0,
			o0 => Or216880_o0
		);
		And216900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216880_o0,
			i1 => i19,
			o0 => And216900_o0
		);
		Or216920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216900_o0,
			i1 => Xor216780_o0,
			o0 => Or216920_o0
		);
		And216940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24940_o0,
			i1 => Nor21260_o0,
			o0 => And216940_o0
		);
		And216960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216940_o0,
			i1 => Or216920_o0,
			o0 => And216960_o0
		);
		Or216980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216960_o0,
			i1 => And216760_o0,
			o0 => Or216980_o0
		);
		And217000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or216980_o0,
			i1 => Not1280_o0,
			o0 => And217000_o0
		);
		Or217020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210020_o0,
			i1 => i19,
			o0 => Or217020_o0
		);
		And217040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217020_o0,
			i1 => i17,
			o0 => And217040_o0
		);
		Or217060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217040_o0,
			i1 => Nor214120_o0,
			o0 => Or217060_o0
		);
		Or217080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or217060_o0,
			i1 => i18,
			o0 => Or217080_o0
		);
		And217100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216700_o0,
			i1 => And2640_o0,
			o0 => And217100_o0
		);
		And217120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217100_o0,
			i1 => Or217080_o0,
			o0 => And217120_o0
		);
		Or217140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217120_o0,
			i1 => And217000_o0,
			o0 => Or217140_o0
		);
		And217160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => Not100_o0,
			o0 => And217160_o0
		);
		And217180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217160_o0,
			i1 => Not2080_o0,
			o0 => And217180_o0
		);
		And217200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217180_o0,
			i1 => Or217140_o0,
			o0 => And217200_o0
		);
		Or217220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217200_o0,
			i1 => And216480_o0,
			o0 => Or217220_o0
		);
		And217240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217220_o0,
			i1 => Not80_o0,
			o0 => And217240_o0
		);
		And217260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22800_o0,
			i1 => Xor2960_o0,
			o0 => And217260_o0
		);
		And217280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => Not620_o0,
			o0 => And217280_o0
		);
		Or217300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217280_o0,
			i1 => And217260_o0,
			o0 => Or217300_o0
		);
		And217320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217300_o0,
			i1 => i18,
			o0 => And217320_o0
		);
		And217340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => i17,
			o0 => And217340_o0
		);
		And217360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217340_o0,
			i1 => Nor21840_o0,
			o0 => And217360_o0
		);
		Or217380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217360_o0,
			i1 => And217320_o0,
			o0 => Or217380_o0
		);
		And217400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217380_o0,
			i1 => i13,
			o0 => And217400_o0
		);
		Nand217420 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i18,
			o0 => Nand217420_o0
		);
		And217440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand217420_o0,
			i1 => Not1280_o0,
			o0 => And217440_o0
		);
		And217460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => i16,
			o0 => And217460_o0
		);
		Or217480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217460_o0,
			i1 => And217440_o0,
			o0 => Or217480_o0
		);
		And217500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i13,
			o0 => And217500_o0
		);
		And217520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217500_o0,
			i1 => Or217480_o0,
			o0 => And217520_o0
		);
		Or217540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217520_o0,
			i1 => Not2080_o0,
			o0 => Or217540_o0
		);
		Or217560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or217540_o0,
			i1 => And217400_o0,
			o0 => Or217560_o0
		);
		And217580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217560_o0,
			i1 => i12,
			o0 => And217580_o0
		);
		And217600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212900_o0,
			i1 => Nor211040_o0,
			o0 => And217600_o0
		);
		Or217620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217600_o0,
			i1 => i13,
			o0 => Or217620_o0
		);
		And217640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217620_o0,
			i1 => Not180_o0,
			o0 => And217640_o0
		);
		Or217660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217640_o0,
			i1 => And217580_o0,
			o0 => Or217660_o0
		);
		And217680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => i14,
			o0 => And217680_o0
		);
		And217700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217680_o0,
			i1 => Nor25100_o0,
			o0 => And217700_o0
		);
		And217720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217700_o0,
			i1 => Or217660_o0,
			o0 => And217720_o0
		);
		Or217740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217720_o0,
			i1 => And217240_o0,
			o0 => Or217740_o0
		);
		And217760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217740_o0,
			i1 => Not140_o0,
			o0 => And217760_o0
		);
		And217780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i23,
			i1 => i22,
			o0 => And217780_o0
		);
		And217800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217780_o0,
			i1 => Not7120_o0,
			o0 => And217800_o0
		);
		Or217820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217800_o0,
			i1 => And210740_o0,
			o0 => Or217820_o0
		);
		Xor217840 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => Not160_o0,
			o0 => Xor217840_o0
		);
		And217860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor217840_o0,
			i1 => Or217820_o0,
			o0 => And217860_o0
		);
		Nand217880 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i25,
			i1 => i23,
			o0 => Nand217880_o0
		);
		Nor217900 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i4,
			o0 => Nor217900_o0
		);
		And217920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => i22,
			o0 => And217920_o0
		);
		And217940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217920_o0,
			i1 => Nor217900_o0,
			o0 => And217940_o0
		);
		And217960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217940_o0,
			i1 => Nand217880_o0,
			o0 => And217960_o0
		);
		Or217980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217960_o0,
			i1 => And217860_o0,
			o0 => Or217980_o0
		);
		And218000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217980_o0,
			i1 => Not540_o0,
			o0 => And218000_o0
		);
		Xor218020 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i24,
			o0 => Xor218020_o0
		);
		Nor218040 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor218020_o0,
			i1 => i23,
			o0 => Nor218040_o0
		);
		Or218060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i25,
			o0 => Or218060_o0
		);
		And218080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218060_o0,
			i1 => i24,
			o0 => And218080_o0
		);
		And218100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218080_o0,
			i1 => i23,
			o0 => And218100_o0
		);
		Or218120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218100_o0,
			i1 => Nor218040_o0,
			o0 => Or218120_o0
		);
		And218140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218120_o0,
			i1 => i22,
			o0 => And218140_o0
		);
		And218160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29640_o0,
			i1 => Not9800_o0,
			o0 => And218160_o0
		);
		Or218180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218160_o0,
			i1 => And218140_o0,
			o0 => Or218180_o0
		);
		And218200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218180_o0,
			i1 => And215860_o0,
			o0 => And218200_o0
		);
		Or218220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218200_o0,
			i1 => And218000_o0,
			o0 => Or218220_o0
		);
		And218240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218220_o0,
			i1 => And29560_o0,
			o0 => And218240_o0
		);
		Nor218260 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i21,
			o0 => Nor218260_o0
		);
		And218280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor218260_o0,
			i1 => i20,
			o0 => And218280_o0
		);
		And218300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218280_o0,
			i1 => And215860_o0,
			o0 => And218300_o0
		);
		Or218320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218300_o0,
			i1 => And218240_o0,
			o0 => Or218320_o0
		);
		And218340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218320_o0,
			i1 => i18,
			o0 => And218340_o0
		);
		And218360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not1080_o0,
			o0 => And218360_o0
		);
		Or218380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218360_o0,
			i1 => And218340_o0,
			o0 => Or218380_o0
		);
		And218400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => Not1500_o0,
			o0 => And218400_o0
		);
		And218420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => And26680_o0,
			o0 => And218420_o0
		);
		And218440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218420_o0,
			i1 => And217160_o0,
			o0 => And218440_o0
		);
		And218460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218440_o0,
			i1 => And218400_o0,
			o0 => And218460_o0
		);
		And218480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218460_o0,
			i1 => Or218380_o0,
			o0 => And218480_o0
		);
		Or218500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218480_o0,
			i1 => And217760_o0,
			o0 => Or218500_o0
		);
		And218520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218500_o0,
			i1 => Not60_o0,
			o0 => And218520_o0
		);
		And218540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or22840_o0,
			i1 => i3,
			o0 => And218540_o0
		);
		And218560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not140_o0,
			o0 => And218560_o0
		);
		And218580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => Not1040_o0,
			o0 => And218580_o0
		);
		And218600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => And218560_o0,
			o0 => And218600_o0
		);
		Or218620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218600_o0,
			i1 => And218540_o0,
			o0 => Or218620_o0
		);
		And218640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218620_o0,
			i1 => i16,
			o0 => And218640_o0
		);
		And218660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21300_o0,
			i1 => Not140_o0,
			o0 => And218660_o0
		);
		And218680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218660_o0,
			i1 => And21240_o0,
			o0 => And218680_o0
		);
		Or218700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218680_o0,
			i1 => And218640_o0,
			o0 => Or218700_o0
		);
		And218720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218700_o0,
			i1 => And23020_o0,
			o0 => And218720_o0
		);
		And218740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => And24140_o0,
			o0 => And218740_o0
		);
		And218760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218740_o0,
			i1 => And21960_o0,
			o0 => And218760_o0
		);
		Or218780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218760_o0,
			i1 => And218720_o0,
			o0 => Or218780_o0
		);
		And218800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not80_o0,
			o0 => And218800_o0
		);
		And218820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218800_o0,
			i1 => And23180_o0,
			o0 => And218820_o0
		);
		And218840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218820_o0,
			i1 => Or218780_o0,
			o0 => And218840_o0
		);
		Or218860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218840_o0,
			i1 => And218520_o0,
			o0 => Or218860_o0
		);
		And218880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or218860_o0,
			i1 => Not120_o0,
			o0 => And218880_o0
		);
		And218900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210600_o0,
			i1 => Not540_o0,
			o0 => And218900_o0
		);
		And218920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210540_o0,
			i1 => i5,
			o0 => And218920_o0
		);
		Or218940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218920_o0,
			i1 => And218900_o0,
			o0 => Or218940_o0
		);
		And218960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => i27,
			o0 => And218960_o0
		);
		And218980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => And21940_o0,
			o0 => And218980_o0
		);
		And219000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218980_o0,
			i1 => And23080_o0,
			o0 => And219000_o0
		);
		And219020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219000_o0,
			i1 => And218960_o0,
			o0 => And219020_o0
		);
		And219040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219020_o0,
			i1 => Or218940_o0,
			o0 => And219040_o0
		);
		And219060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not140_o0,
			i1 => i2,
			o0 => And219060_o0
		);
		And219080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219060_o0,
			i1 => Not160_o0,
			o0 => And219080_o0
		);
		And219100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219080_o0,
			i1 => Nor23600_o0,
			o0 => And219100_o0
		);
		And219120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219100_o0,
			i1 => And219040_o0,
			o0 => And219120_o0
		);
		Or219140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219120_o0,
			i1 => And218880_o0,
			o0 => Or219140_o0
		);
		And219160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219140_o0,
			i1 => And23360_o0,
			o0 => And219160_o0
		);
		Or219180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => i16,
			o0 => Or219180_o0
		);
		Or219200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or219180_o0,
			i1 => Not2080_o0,
			o0 => Or219200_o0
		);
		And219220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219200_o0,
			i1 => Not1040_o0,
			o0 => And219220_o0
		);
		Or219240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not2080_o0,
			o0 => Or219240_o0
		);
		And219260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219240_o0,
			i1 => i17,
			o0 => And219260_o0
		);
		Or219280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219260_o0,
			i1 => And219220_o0,
			o0 => Or219280_o0
		);
		And219300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219280_o0,
			i1 => i18,
			o0 => And219300_o0
		);
		Or219320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210420_o0,
			i1 => Not2080_o0,
			o0 => Or219320_o0
		);
		And219340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219320_o0,
			i1 => Not1080_o0,
			o0 => And219340_o0
		);
		Or219360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219340_o0,
			i1 => And219300_o0,
			o0 => Or219360_o0
		);
		And219380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219360_o0,
			i1 => i15,
			o0 => And219380_o0
		);
		Or219400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219380_o0,
			i1 => Nor211040_o0,
			o0 => Or219400_o0
		);
		And219420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219400_o0,
			i1 => Not80_o0,
			o0 => And219420_o0
		);
		And219440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219420_o0,
			i1 => Not540_o0,
			o0 => And219440_o0
		);
		Or219460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i15,
			o0 => Or219460_o0
		);
		Or219480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or219460_o0,
			i1 => And217280_o0,
			o0 => Or219480_o0
		);
		And219500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not2080_o0,
			i1 => i5,
			o0 => And219500_o0
		);
		And219520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219500_o0,
			i1 => i14,
			o0 => And219520_o0
		);
		And219540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219520_o0,
			i1 => Or219480_o0,
			o0 => And219540_o0
		);
		Or219560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219540_o0,
			i1 => And219440_o0,
			o0 => Or219560_o0
		);
		And219580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219560_o0,
			i1 => Not180_o0,
			o0 => And219580_o0
		);
		And219600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i13,
			o0 => And219600_o0
		);
		And219620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not80_o0,
			o0 => And219620_o0
		);
		And219640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219620_o0,
			i1 => Not2080_o0,
			o0 => And219640_o0
		);
		Or219660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219640_o0,
			i1 => And219600_o0,
			o0 => Or219660_o0
		);
		And219680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219660_o0,
			i1 => i17,
			o0 => And219680_o0
		);
		And219700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => And21060_o0,
			o0 => And219700_o0
		);
		Or219720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219700_o0,
			i1 => And219680_o0,
			o0 => Or219720_o0
		);
		And219740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219720_o0,
			i1 => i15,
			o0 => And219740_o0
		);
		And219760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => And210440_o0,
			o0 => And219760_o0
		);
		And219780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => i13,
			o0 => And219780_o0
		);
		And219800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => i16,
			o0 => And219800_o0
		);
		And219820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219800_o0,
			i1 => And219780_o0,
			o0 => And219820_o0
		);
		Or219840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219820_o0,
			i1 => And219760_o0,
			o0 => Or219840_o0
		);
		Or219860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or219840_o0,
			i1 => And219740_o0,
			o0 => Or219860_o0
		);
		And219880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219860_o0,
			i1 => And211020_o0,
			o0 => And219880_o0
		);
		And219900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not80_o0,
			o0 => And219900_o0
		);
		And219920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => Not2080_o0,
			o0 => And219920_o0
		);
		And219940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => Not1280_o0,
			o0 => And219940_o0
		);
		And219960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219940_o0,
			i1 => And219920_o0,
			o0 => And219960_o0
		);
		And219980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219780_o0,
			i1 => And2320_o0,
			o0 => And219980_o0
		);
		Or220000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219980_o0,
			i1 => And219960_o0,
			o0 => Or220000_o0
		);
		And220020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220000_o0,
			i1 => i5,
			o0 => And220020_o0
		);
		And220040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => Not1080_o0,
			o0 => And220040_o0
		);
		Nor220060 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => i5,
			o0 => Nor220060_o0
		);
		And220080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216820_o0,
			i1 => Nor24920_o0,
			o0 => And220080_o0
		);
		And220100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220080_o0,
			i1 => Nor220060_o0,
			o0 => And220100_o0
		);
		And220120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220100_o0,
			i1 => And220040_o0,
			o0 => And220120_o0
		);
		Or220140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220120_o0,
			i1 => And220020_o0,
			o0 => Or220140_o0
		);
		And220160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220140_o0,
			i1 => i19,
			o0 => And220160_o0
		);
		And220180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => Nor21220_o0,
			o0 => And220180_o0
		);
		And220200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => Nor22900_o0,
			o0 => And220200_o0
		);
		And220220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220200_o0,
			i1 => Nor220060_o0,
			o0 => And220220_o0
		);
		And220240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220220_o0,
			i1 => And220180_o0,
			o0 => And220240_o0
		);
		Or220260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220240_o0,
			i1 => And220160_o0,
			o0 => Or220260_o0
		);
		And220280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220260_o0,
			i1 => i12,
			o0 => And220280_o0
		);
		Or220300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220280_o0,
			i1 => And219880_o0,
			o0 => Or220300_o0
		);
		Or220320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or220300_o0,
			i1 => And219580_o0,
			o0 => Or220320_o0
		);
		Nor220340 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i9,
			i1 => i4,
			o0 => Nor220340_o0
		);
		And220360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor220340_o0,
			i1 => Nor21140_o0,
			o0 => And220360_o0
		);
		And220380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220360_o0,
			i1 => Nor23600_o0,
			o0 => And220380_o0
		);
		And220400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220380_o0,
			i1 => And213240_o0,
			o0 => And220400_o0
		);
		And220420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220400_o0,
			i1 => Or220320_o0,
			o0 => And220420_o0
		);
		And220440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			i1 => i10,
			o0 => And220440_o0
		);
		And220460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220440_o0,
			i1 => i9,
			o0 => And220460_o0
		);
		Or220480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220460_o0,
			i1 => And220420_o0,
			o0 => Or220480_o0
		);
		And220500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220480_o0,
			i1 => Not12100_o0,
			o0 => And220500_o0
		);
		Not20520 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i9,
			o0 => Not20520_o0
		);
		And220540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not3300_o0,
			i1 => i8,
			o0 => And220540_o0
		);
		And220560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220540_o0,
			i1 => Nor21260_o0,
			o0 => And220560_o0
		);
		And220580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220560_o0,
			i1 => And28160_o0,
			o0 => And220580_o0
		);
		And220600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => Not12100_o0,
			o0 => And220600_o0
		);
		Or220620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220600_o0,
			i1 => And220580_o0,
			o0 => Or220620_o0
		);
		And220640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220620_o0,
			i1 => Not20520_o0,
			o0 => And220640_o0
		);
		And220660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12120_o0,
			i1 => i9,
			o0 => And220660_o0
		);
		And220680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220660_o0,
			i1 => Not12100_o0,
			o0 => And220680_o0
		);
		Or220700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => o71,
			i1 => And220640_o0,
			o0 => Or220700_o0
		);
		Or220720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or220700_o0,
			i1 => And220500_o0,
			o0 => Or220720_o0
		);
		And220740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => i9,
			o0 => And220740_o0
		);
		Not20760 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			o0 => Not20760_o0
		);
		Or220780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And210440_o0,
			i1 => And23780_o0,
			o0 => Or220780_o0
		);
		And220800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220780_o0,
			i1 => Not20760_o0,
			o0 => And220800_o0
		);
		And220820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212280_o0,
			i1 => And22800_o0,
			o0 => And220820_o0
		);
		Or220840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220820_o0,
			i1 => And22300_o0,
			o0 => Or220840_o0
		);
		And220860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220840_o0,
			i1 => Not1280_o0,
			o0 => And220860_o0
		);
		Or220880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220860_o0,
			i1 => And220800_o0,
			o0 => Or220880_o0
		);
		And220900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220880_o0,
			i1 => Not1080_o0,
			o0 => And220900_o0
		);
		Or220920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			i1 => i20,
			o0 => Or220920_o0
		);
		And220940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220920_o0,
			i1 => i18,
			o0 => And220940_o0
		);
		And220960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220940_o0,
			i1 => And29520_o0,
			o0 => And220960_o0
		);
		Or220980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And220960_o0,
			i1 => And220900_o0,
			o0 => Or220980_o0
		);
		And221000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220980_o0,
			i1 => And2560_o0,
			o0 => And221000_o0
		);
		Xor221020 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			i1 => i20,
			o0 => Xor221020_o0
		);
		Or221040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Xor221020_o0,
			i1 => Not1080_o0,
			o0 => Or221040_o0
		);
		And221060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221040_o0,
			i1 => And29520_o0,
			o0 => And221060_o0
		);
		And221080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221060_o0,
			i1 => i5,
			o0 => And221080_o0
		);
		Or221100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221080_o0,
			i1 => And221000_o0,
			o0 => Or221100_o0
		);
		And221120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221100_o0,
			i1 => Not160_o0,
			o0 => And221120_o0
		);
		And221140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221060_o0,
			i1 => i4,
			o0 => And221140_o0
		);
		Or221160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221140_o0,
			i1 => And221120_o0,
			o0 => Or221160_o0
		);
		And221180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221160_o0,
			i1 => Not140_o0,
			o0 => And221180_o0
		);
		Or221200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => Not7120_o0,
			o0 => Or221200_o0
		);
		And221220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221200_o0,
			i1 => Nand210560_o0,
			o0 => And221220_o0
		);
		And221240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => Not7120_o0,
			o0 => And221240_o0
		);
		Or221260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221240_o0,
			i1 => And218080_o0,
			o0 => Or221260_o0
		);
		And221280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221260_o0,
			i1 => And217780_o0,
			o0 => And221280_o0
		);
		Or221300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221280_o0,
			i1 => And221220_o0,
			o0 => Or221300_o0
		);
		And221320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221300_o0,
			i1 => Not540_o0,
			o0 => And221320_o0
		);
		Nand221340 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => i22,
			o0 => Nand221340_o0
		);
		And221360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i5,
			o0 => And221360_o0
		);
		And221380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221360_o0,
			i1 => Nand221340_o0,
			o0 => And221380_o0
		);
		Or221400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221380_o0,
			i1 => And221320_o0,
			o0 => Or221400_o0
		);
		And221420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221400_o0,
			i1 => Not160_o0,
			o0 => And221420_o0
		);
		And221440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210560_o0,
			i1 => i27,
			o0 => And221440_o0
		);
		And221460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221440_o0,
			i1 => Not7120_o0,
			o0 => And221460_o0
		);
		And221480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221460_o0,
			i1 => i4,
			o0 => And221480_o0
		);
		Or221500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221480_o0,
			i1 => And221420_o0,
			o0 => Or221500_o0
		);
		And221520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221500_o0,
			i1 => And29560_o0,
			o0 => And221520_o0
		);
		Or221540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => i27,
			o0 => Or221540_o0
		);
		And221560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221540_o0,
			i1 => And210540_o0,
			o0 => And221560_o0
		);
		Or221580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221560_o0,
			i1 => And221520_o0,
			o0 => Or221580_o0
		);
		And221600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => i18,
			o0 => And221600_o0
		);
		And221620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221600_o0,
			i1 => And26680_o0,
			o0 => And221620_o0
		);
		And221640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221620_o0,
			i1 => Or221580_o0,
			o0 => And221640_o0
		);
		Or221660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221640_o0,
			i1 => And221180_o0,
			o0 => Or221660_o0
		);
		And221680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221660_o0,
			i1 => Not1500_o0,
			o0 => And221680_o0
		);
		And221700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i15,
			o0 => And221700_o0
		);
		And221720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => Not1080_o0,
			o0 => And221720_o0
		);
		And221740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221720_o0,
			i1 => And22300_o0,
			o0 => And221740_o0
		);
		Or221760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221740_o0,
			i1 => And221700_o0,
			o0 => Or221760_o0
		);
		And221780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221760_o0,
			i1 => And2560_o0,
			o0 => And221780_o0
		);
		And221800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => And28460_o0,
			o0 => And221800_o0
		);
		Or221820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221800_o0,
			i1 => And221780_o0,
			o0 => Or221820_o0
		);
		And221840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221820_o0,
			i1 => Not160_o0,
			o0 => And221840_o0
		);
		And221860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214860_o0,
			i1 => i15,
			o0 => And221860_o0
		);
		And221880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221860_o0,
			i1 => And212880_o0,
			o0 => And221880_o0
		);
		Or221900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221880_o0,
			i1 => And221840_o0,
			o0 => Or221900_o0
		);
		Nor221920 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i3,
			o0 => Nor221920_o0
		);
		And221940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor221920_o0,
			i1 => i19,
			o0 => And221940_o0
		);
		And221960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221940_o0,
			i1 => Or221900_o0,
			o0 => And221960_o0
		);
		Or221980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And221960_o0,
			i1 => And221680_o0,
			o0 => Or221980_o0
		);
		And222000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221980_o0,
			i1 => And23080_o0,
			o0 => And222000_o0
		);
		And222020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215820_o0,
			i1 => Not620_o0,
			o0 => And222020_o0
		);
		And222040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215880_o0,
			i1 => i15,
			o0 => And222040_o0
		);
		Or222060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222040_o0,
			i1 => And222020_o0,
			o0 => Or222060_o0
		);
		And222080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210400_o0,
			i1 => i18,
			o0 => And222080_o0
		);
		And222100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222080_o0,
			i1 => Or222060_o0,
			o0 => And222100_o0
		);
		And222120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not1500_o0,
			o0 => And222120_o0
		);
		And222140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222120_o0,
			i1 => Not1080_o0,
			o0 => And222140_o0
		);
		And222160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => Not540_o0,
			o0 => And222160_o0
		);
		And222180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222160_o0,
			i1 => And222140_o0,
			o0 => And222180_o0
		);
		Or222200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222180_o0,
			i1 => And222100_o0,
			o0 => Or222200_o0
		);
		And222220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222200_o0,
			i1 => Not160_o0,
			o0 => And222220_o0
		);
		And222240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i4,
			o0 => And222240_o0
		);
		And222260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222240_o0,
			i1 => Or222060_o0,
			o0 => And222260_o0
		);
		Or222280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222260_o0,
			i1 => And222220_o0,
			o0 => Or222280_o0
		);
		And222300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222280_o0,
			i1 => Not140_o0,
			o0 => And222300_o0
		);
		And222320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2240_o0,
			i1 => i16,
			o0 => And222320_o0
		);
		And222340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222320_o0,
			i1 => And26680_o0,
			o0 => And222340_o0
		);
		Or222360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222340_o0,
			i1 => And222300_o0,
			o0 => Or222360_o0
		);
		And222380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => i17,
			o0 => And222380_o0
		);
		And222400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222380_o0,
			i1 => Or222360_o0,
			o0 => And222400_o0
		);
		Or222420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222400_o0,
			i1 => And222000_o0,
			o0 => Or222420_o0
		);
		And222440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222420_o0,
			i1 => Not100_o0,
			o0 => And222440_o0
		);
		And222460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25020_o0,
			i1 => And21000_o0,
			o0 => And222460_o0
		);
		And222480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => Not140_o0,
			o0 => And222480_o0
		);
		And222500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222480_o0,
			i1 => And2260_o0,
			o0 => And222500_o0
		);
		And222520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28460_o0,
			i1 => Nor22600_o0,
			o0 => And222520_o0
		);
		And222540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222520_o0,
			i1 => And22920_o0,
			o0 => And222540_o0
		);
		Or222560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222540_o0,
			i1 => And222500_o0,
			o0 => Or222560_o0
		);
		Or222580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or222560_o0,
			i1 => And222460_o0,
			o0 => Or222580_o0
		);
		Or222600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or222580_o0,
			i1 => And27400_o0,
			o0 => Or222600_o0
		);
		And222620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222600_o0,
			i1 => And211600_o0,
			o0 => And222620_o0
		);
		Or222640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222620_o0,
			i1 => And222440_o0,
			o0 => Or222640_o0
		);
		And222660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222640_o0,
			i1 => Not120_o0,
			o0 => And222660_o0
		);
		And222680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or21020_o0,
			i1 => i1,
			o0 => And222680_o0
		);
		And222700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => Not100_o0,
			o0 => And222700_o0
		);
		And222720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222700_o0,
			i1 => And2260_o0,
			o0 => And222720_o0
		);
		Or222740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222720_o0,
			i1 => And222680_o0,
			o0 => Or222740_o0
		);
		And222760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222740_o0,
			i1 => And23020_o0,
			o0 => And222760_o0
		);
		And222780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => Nor22600_o0,
			o0 => And222780_o0
		);
		And222800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => Not540_o0,
			o0 => And222800_o0
		);
		And222820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => Not10520_o0,
			o0 => And222820_o0
		);
		And222840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222820_o0,
			i1 => And222800_o0,
			o0 => And222840_o0
		);
		And222860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222840_o0,
			i1 => And222780_o0,
			o0 => And222860_o0
		);
		Nor222880 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i1,
			o0 => Nor222880_o0
		);
		And222900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor222880_o0,
			i1 => i20,
			o0 => And222900_o0
		);
		And222920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222900_o0,
			i1 => And219940_o0,
			o0 => And222920_o0
		);
		And222940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222920_o0,
			i1 => And222860_o0,
			o0 => And222940_o0
		);
		Or222960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222940_o0,
			i1 => And222760_o0,
			o0 => Or222960_o0
		);
		And222980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or222960_o0,
			i1 => i2,
			o0 => And222980_o0
		);
		Or223000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222980_o0,
			i1 => And222660_o0,
			o0 => Or223000_o0
		);
		And223020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223000_o0,
			i1 => Not80_o0,
			o0 => And223020_o0
		);
		Or223040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or210400_o0,
			i1 => i4,
			o0 => Or223040_o0
		);
		And223060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223040_o0,
			i1 => And23520_o0,
			o0 => And223060_o0
		);
		And223080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not2080_o0,
			o0 => And223080_o0
		);
		And223100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223080_o0,
			i1 => And24040_o0,
			o0 => And223100_o0
		);
		Or223120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223100_o0,
			i1 => And223060_o0,
			o0 => Or223120_o0
		);
		And223140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223120_o0,
			i1 => Not1080_o0,
			o0 => And223140_o0
		);
		And223160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor220060_o0,
			i1 => Not160_o0,
			o0 => And223160_o0
		);
		And223180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223160_o0,
			i1 => And24200_o0,
			o0 => And223180_o0
		);
		Or223200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223180_o0,
			i1 => And223140_o0,
			o0 => Or223200_o0
		);
		And223220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223200_o0,
			i1 => Not1040_o0,
			o0 => And223220_o0
		);
		And223240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i17,
			o0 => And223240_o0
		);
		And223260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => Not2080_o0,
			o0 => And223260_o0
		);
		And223280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223260_o0,
			i1 => Nor21260_o0,
			o0 => And223280_o0
		);
		And223300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223280_o0,
			i1 => And223240_o0,
			o0 => And223300_o0
		);
		Or223320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223300_o0,
			i1 => And223220_o0,
			o0 => Or223320_o0
		);
		And223340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223320_o0,
			i1 => i15,
			o0 => And223340_o0
		);
		Or223360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not1080_o0,
			i1 => i17,
			o0 => Or223360_o0
		);
		And223380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not620_o0,
			o0 => And223380_o0
		);
		And223400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223380_o0,
			i1 => And223260_o0,
			o0 => And223400_o0
		);
		And223420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223400_o0,
			i1 => Nor21260_o0,
			o0 => And223420_o0
		);
		And223440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223420_o0,
			i1 => Or223360_o0,
			o0 => And223440_o0
		);
		Or223460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223440_o0,
			i1 => And223340_o0,
			o0 => Or223460_o0
		);
		And223480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223460_o0,
			i1 => Not180_o0,
			o0 => And223480_o0
		);
		And223500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => And28060_o0,
			o0 => And223500_o0
		);
		And223520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223240_o0,
			i1 => Nor21260_o0,
			o0 => And223520_o0
		);
		And223540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223520_o0,
			i1 => And223500_o0,
			o0 => And223540_o0
		);
		Or223560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223540_o0,
			i1 => And223480_o0,
			o0 => Or223560_o0
		);
		And223580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223560_o0,
			i1 => Not140_o0,
			o0 => And223580_o0
		);
		And223600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Not80_o0,
			o0 => And223600_o0
		);
		And223620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223600_o0,
			i1 => And2600_o0,
			o0 => And223620_o0
		);
		And223640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223620_o0,
			i1 => i3,
			o0 => And223640_o0
		);
		Or223660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223640_o0,
			i1 => And223580_o0,
			o0 => Or223660_o0
		);
		And223680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223660_o0,
			i1 => Not120_o0,
			o0 => And223680_o0
		);
		And223700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223620_o0,
			i1 => i2,
			o0 => And223700_o0
		);
		Or223720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223700_o0,
			i1 => And223680_o0,
			o0 => Or223720_o0
		);
		And223740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223720_o0,
			i1 => Not100_o0,
			o0 => And223740_o0
		);
		And223760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223040_o0,
			i1 => And210100_o0,
			o0 => And223760_o0
		);
		Nand223780 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => i37,
			o0 => Nand223780_o0
		);
		And223800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216700_o0,
			i1 => And212880_o0,
			o0 => And223800_o0
		);
		And223820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223800_o0,
			i1 => Nand223780_o0,
			o0 => And223820_o0
		);
		Or223840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223820_o0,
			i1 => And223760_o0,
			o0 => Or223840_o0
		);
		And223860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Not1280_o0,
			o0 => And223860_o0
		);
		And223880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223860_o0,
			i1 => Or223840_o0,
			o0 => And223880_o0
		);
		And223900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28480_o0,
			i1 => And27940_o0,
			o0 => And223900_o0
		);
		Or223920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And223900_o0,
			i1 => And223880_o0,
			o0 => Or223920_o0
		);
		And223940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223920_o0,
			i1 => And219900_o0,
			o0 => And223940_o0
		);
		Or223960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i17,
			o0 => Or223960_o0
		);
		And223980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223960_o0,
			i1 => And28120_o0,
			o0 => And223980_o0
		);
		Nor224000 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => i12,
			o0 => Nor224000_o0
		);
		And224020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor224000_o0,
			i1 => And212880_o0,
			o0 => And224020_o0
		);
		Or224040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224020_o0,
			i1 => And223980_o0,
			o0 => Or224040_o0
		);
		And224060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => And28480_o0,
			o0 => And224060_o0
		);
		And224080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224060_o0,
			i1 => Nor21260_o0,
			o0 => And224080_o0
		);
		And224100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224080_o0,
			i1 => Or224040_o0,
			o0 => And224100_o0
		);
		Or224120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224100_o0,
			i1 => And223940_o0,
			o0 => Or224120_o0
		);
		And224140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or224120_o0,
			i1 => Not140_o0,
			o0 => And224140_o0
		);
		And224160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210100_o0,
			i1 => Not1280_o0,
			o0 => And224160_o0
		);
		And224180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224160_o0,
			i1 => And219900_o0,
			o0 => And224180_o0
		);
		And224200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not160_o0,
			i1 => i3,
			o0 => And224200_o0
		);
		And224220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Not540_o0,
			o0 => And224220_o0
		);
		And224240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224220_o0,
			i1 => And224200_o0,
			o0 => And224240_o0
		);
		And224260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224240_o0,
			i1 => And224180_o0,
			o0 => And224260_o0
		);
		Or224280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224260_o0,
			i1 => And224140_o0,
			o0 => Or224280_o0
		);
		And224300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or224280_o0,
			i1 => Not100_o0,
			o0 => And224300_o0
		);
		And224320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => Not140_o0,
			o0 => And224320_o0
		);
		And224340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224320_o0,
			i1 => And25300_o0,
			o0 => And224340_o0
		);
		And224360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => And24280_o0,
			o0 => And224360_o0
		);
		And224380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224360_o0,
			i1 => And224340_o0,
			o0 => And224380_o0
		);
		And224400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224380_o0,
			i1 => And2320_o0,
			o0 => And224400_o0
		);
		Or224420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224400_o0,
			i1 => And224300_o0,
			o0 => Or224420_o0
		);
		And224440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or224420_o0,
			i1 => Not120_o0,
			o0 => And224440_o0
		);
		And224460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not120_o0,
			i1 => i1,
			o0 => And224460_o0
		);
		And224480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224460_o0,
			i1 => And2600_o0,
			o0 => And224480_o0
		);
		And224500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => Not180_o0,
			o0 => And224500_o0
		);
		And224520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224500_o0,
			i1 => And24860_o0,
			o0 => And224520_o0
		);
		And224540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224520_o0,
			i1 => And224480_o0,
			o0 => And224540_o0
		);
		Not24560 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			o0 => Not24560_o0
		);
		And224580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i19,
			o0 => And224580_o0
		);
		And224600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => Not1080_o0,
			o0 => And224600_o0
		);
		And224620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => And21060_o0,
			o0 => And224620_o0
		);
		And224640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224620_o0,
			i1 => And213180_o0,
			o0 => And224640_o0
		);
		And224660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224640_o0,
			i1 => And224600_o0,
			o0 => And224660_o0
		);
		Or224680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224660_o0,
			i1 => Not24560_o0,
			o0 => Or224680_o0
		);
		And224700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22600_o0,
			i1 => Not540_o0,
			o0 => And224700_o0
		);
		And224720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224700_o0,
			i1 => Nor22060_o0,
			o0 => And224720_o0
		);
		And224740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224720_o0,
			i1 => Or224680_o0,
			o0 => And224740_o0
		);
		Or224760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224740_o0,
			i1 => And224540_o0,
			o0 => Or224760_o0
		);
		Or224780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or224760_o0,
			i1 => And224440_o0,
			o0 => Or224780_o0
		);
		Or224800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or224780_o0,
			i1 => And223740_o0,
			o0 => Or224800_o0
		);
		Or224820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or224800_o0,
			i1 => And223020_o0,
			o0 => Or224820_o0
		);
		And224840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or224820_o0,
			i1 => Not60_o0,
			o0 => And224840_o0
		);
		Or224860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28920_o0,
			i1 => And22860_o0,
			o0 => Or224860_o0
		);
		And224880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223600_o0,
			i1 => And211740_o0,
			o0 => And224880_o0
		);
		And224900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224880_o0,
			i1 => Or224860_o0,
			o0 => And224900_o0
		);
		Or224920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224900_o0,
			i1 => And224840_o0,
			o0 => Or224920_o0
		);
		Or224940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or224920_o0,
			i1 => i36,
			o0 => Or224940_o0
		);
		Not24960 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			o0 => Not24960_o0
		);
		And224980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212700_o0,
			i1 => Not24960_o0,
			o0 => And224980_o0
		);
		And225000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224980_o0,
			i1 => Or224940_o0,
			o0 => And225000_o0
		);
		Or225020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225000_o0,
			i1 => And220740_o0,
			o0 => Or225020_o0
		);
		And225040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225020_o0,
			i1 => Not12100_o0,
			o0 => And225040_o0
		);
		And225060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor224000_o0,
			i1 => Not1080_o0,
			o0 => And225060_o0
		);
		And225080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => And2240_o0,
			o0 => And225080_o0
		);
		Or225100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225080_o0,
			i1 => And225060_o0,
			o0 => Or225100_o0
		);
		And225120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225100_o0,
			i1 => Nor21840_o0,
			o0 => And225120_o0
		);
		And225140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => i15,
			o0 => And225140_o0
		);
		And225160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225140_o0,
			i1 => And215820_o0,
			o0 => And225160_o0
		);
		Or225180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225160_o0,
			i1 => And225120_o0,
			o0 => Or225180_o0
		);
		And225200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225180_o0,
			i1 => Not1040_o0,
			o0 => And225200_o0
		);
		And225220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not620_o0,
			i1 => i13,
			o0 => And225220_o0
		);
		And225240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225220_o0,
			i1 => i12,
			o0 => And225240_o0
		);
		And225260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225240_o0,
			i1 => And21960_o0,
			o0 => And225260_o0
		);
		Or225280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225260_o0,
			i1 => And225200_o0,
			o0 => Or225280_o0
		);
		And225300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225280_o0,
			i1 => i14,
			o0 => And225300_o0
		);
		And225320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => i13,
			o0 => And225320_o0
		);
		And225340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => Nor211040_o0,
			o0 => And225340_o0
		);
		Or225360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225340_o0,
			i1 => And225320_o0,
			o0 => Or225360_o0
		);
		And225380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213900_o0,
			i1 => i16,
			o0 => And225380_o0
		);
		And225400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225380_o0,
			i1 => Or225360_o0,
			o0 => And225400_o0
		);
		Or225420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225400_o0,
			i1 => And225300_o0,
			o0 => Or225420_o0
		);
		And225440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225420_o0,
			i1 => And213300_o0,
			o0 => And225440_o0
		);
		And225460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2240_o0,
			i1 => Not1040_o0,
			o0 => And225460_o0
		);
		Or225480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225460_o0,
			i1 => And21820_o0,
			o0 => Or225480_o0
		);
		And225500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225480_o0,
			i1 => And28120_o0,
			o0 => And225500_o0
		);
		And225520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor224000_o0,
			i1 => Nor2220_o0,
			o0 => And225520_o0
		);
		Or225540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225520_o0,
			i1 => And225500_o0,
			o0 => Or225540_o0
		);
		And225560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225540_o0,
			i1 => i14,
			o0 => And225560_o0
		);
		And225580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214400_o0,
			i1 => And21100_o0,
			o0 => And225580_o0
		);
		And225600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216820_o0,
			i1 => And23080_o0,
			o0 => And225600_o0
		);
		And225620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225600_o0,
			i1 => And225580_o0,
			o0 => And225620_o0
		);
		Or225640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225620_o0,
			i1 => And225560_o0,
			o0 => Or225640_o0
		);
		And225660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225640_o0,
			i1 => Not620_o0,
			o0 => And225660_o0
		);
		And225680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i13,
			o0 => And225680_o0
		);
		And225700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225680_o0,
			i1 => Not180_o0,
			o0 => And225700_o0
		);
		And225720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Nor21220_o0,
			o0 => And225720_o0
		);
		Or225740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225720_o0,
			i1 => And225700_o0,
			o0 => Or225740_o0
		);
		And225760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i37,
			i1 => Not1040_o0,
			o0 => And225760_o0
		);
		And225780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225760_o0,
			i1 => Nor212260_o0,
			o0 => And225780_o0
		);
		And225800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225780_o0,
			i1 => And219900_o0,
			o0 => And225800_o0
		);
		And225820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225800_o0,
			i1 => Or225740_o0,
			o0 => And225820_o0
		);
		Or225840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225820_o0,
			i1 => And225660_o0,
			o0 => Or225840_o0
		);
		Nor225860 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i11,
			o0 => Nor225860_o0
		);
		And225880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor225860_o0,
			i1 => i40,
			o0 => And225880_o0
		);
		And225900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225880_o0,
			i1 => Nor214960_o0,
			o0 => And225900_o0
		);
		And225920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225900_o0,
			i1 => Or225840_o0,
			o0 => And225920_o0
		);
		Or225940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And225920_o0,
			i1 => i8,
			o0 => Or225940_o0
		);
		And225960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or225940_o0,
			i1 => Not140_o0,
			o0 => And225960_o0
		);
		And225980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => And21940_o0,
			o0 => And225980_o0
		);
		And226000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225980_o0,
			i1 => Nand217420_o0,
			o0 => And226000_o0
		);
		Nor226020 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i11,
			o0 => Nor226020_o0
		);
		And226040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor226020_o0,
			i1 => i13,
			o0 => And226040_o0
		);
		And226060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226040_o0,
			i1 => Nor214960_o0,
			o0 => And226060_o0
		);
		And226080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226060_o0,
			i1 => And226000_o0,
			o0 => And226080_o0
		);
		And226100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226080_o0,
			i1 => i3,
			o0 => And226100_o0
		);
		Or226120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226100_o0,
			i1 => And225960_o0,
			o0 => Or226120_o0
		);
		Nor226140 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i2,
			o0 => Nor226140_o0
		);
		Nor226160 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i5,
			o0 => Nor226160_o0
		);
		And226180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor226160_o0,
			i1 => Nor226140_o0,
			o0 => And226180_o0
		);
		And226200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226180_o0,
			i1 => Nor23600_o0,
			o0 => And226200_o0
		);
		And226220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226200_o0,
			i1 => Or226120_o0,
			o0 => And226220_o0
		);
		Or226240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226220_o0,
			i1 => And220600_o0,
			o0 => Or226240_o0
		);
		And226260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226240_o0,
			i1 => Not20520_o0,
			o0 => And226260_o0
		);
		And226280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212160_o0,
			i1 => Not12100_o0,
			o0 => And226280_o0
		);
		Or226300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226280_o0,
			i1 => And226260_o0,
			o0 => Or226300_o0
		);
		And226320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => Not2080_o0,
			o0 => And226320_o0
		);
		And226340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => Not1280_o0,
			o0 => And226340_o0
		);
		And226360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226340_o0,
			i1 => And226320_o0,
			o0 => And226360_o0
		);
		Or226380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226360_o0,
			i1 => And219420_o0,
			o0 => Or226380_o0
		);
		And226400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226380_o0,
			i1 => Not180_o0,
			o0 => And226400_o0
		);
		And226420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29940_o0,
			i1 => And22400_o0,
			o0 => And226420_o0
		);
		And226440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => And21520_o0,
			o0 => And226440_o0
		);
		Or226460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226440_o0,
			i1 => And226420_o0,
			o0 => Or226460_o0
		);
		And226480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226460_o0,
			i1 => And219600_o0,
			o0 => And226480_o0
		);
		Nor226500 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i19,
			o0 => Nor226500_o0
		);
		And226520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor226500_o0,
			i1 => And22800_o0,
			o0 => And226520_o0
		);
		And226540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i37,
			i1 => i19,
			o0 => And226540_o0
		);
		And226560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226540_o0,
			i1 => And22300_o0,
			o0 => And226560_o0
		);
		Or226580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226560_o0,
			i1 => And226520_o0,
			o0 => Or226580_o0
		);
		And226600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226580_o0,
			i1 => Not16800_o0,
			o0 => And226600_o0
		);
		And226620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226600_o0,
			i1 => Not1280_o0,
			o0 => And226620_o0
		);
		And226640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29940_o0,
			i1 => And2640_o0,
			o0 => And226640_o0
		);
		Or226660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226640_o0,
			i1 => And226620_o0,
			o0 => Or226660_o0
		);
		And226680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226660_o0,
			i1 => Nor29260_o0,
			o0 => And226680_o0
		);
		Or226700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226680_o0,
			i1 => And226480_o0,
			o0 => Or226700_o0
		);
		And226720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226700_o0,
			i1 => Not1080_o0,
			o0 => And226720_o0
		);
		Xor226740 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not620_o0,
			o0 => Xor226740_o0
		);
		And226760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213700_o0,
			i1 => And29940_o0,
			o0 => And226760_o0
		);
		And226780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226760_o0,
			i1 => Xor226740_o0,
			o0 => And226780_o0
		);
		And226800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22400_o0,
			i1 => Not80_o0,
			o0 => And226800_o0
		);
		Or226820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226800_o0,
			i1 => And226780_o0,
			o0 => Or226820_o0
		);
		And226840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226820_o0,
			i1 => i13,
			o0 => And226840_o0
		);
		Or226860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226840_o0,
			i1 => And226720_o0,
			o0 => Or226860_o0
		);
		And226880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226860_o0,
			i1 => i12,
			o0 => And226880_o0
		);
		Or226900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226880_o0,
			i1 => And226400_o0,
			o0 => Or226900_o0
		);
		And226920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not24960_o0,
			o0 => And226920_o0
		);
		And226940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226920_o0,
			i1 => Nor214960_o0,
			o0 => And226940_o0
		);
		And226960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226940_o0,
			i1 => Or226900_o0,
			o0 => And226960_o0
		);
		Or226980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226960_o0,
			i1 => i8,
			o0 => Or226980_o0
		);
		And227000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or226980_o0,
			i1 => Not540_o0,
			o0 => And227000_o0
		);
		And227020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219460_o0,
			i1 => i14,
			o0 => And227020_o0
		);
		And227040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227020_o0,
			i1 => Not180_o0,
			o0 => And227040_o0
		);
		And227060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213900_o0,
			i1 => And22400_o0,
			o0 => And227060_o0
		);
		Or227080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227060_o0,
			i1 => And227040_o0,
			o0 => Or227080_o0
		);
		And227100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => Not180_o0,
			o0 => And227100_o0
		);
		And227120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227100_o0,
			i1 => And217280_o0,
			o0 => And227120_o0
		);
		Or227140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227120_o0,
			i1 => Or227080_o0,
			o0 => Or227140_o0
		);
		And227160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227140_o0,
			i1 => Not2080_o0,
			o0 => And227160_o0
		);
		And227180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i12,
			o0 => And227180_o0
		);
		And227200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227180_o0,
			i1 => Or220000_o0,
			o0 => And227200_o0
		);
		And227220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219460_o0,
			i1 => i17,
			o0 => And227220_o0
		);
		And227240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => i14,
			o0 => And227240_o0
		);
		And227260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227240_o0,
			i1 => And227220_o0,
			o0 => And227260_o0
		);
		And227280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => And2640_o0,
			o0 => And227280_o0
		);
		And227300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => i12,
			o0 => And227300_o0
		);
		And227320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227300_o0,
			i1 => And227280_o0,
			o0 => And227320_o0
		);
		Or227340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227320_o0,
			i1 => And227260_o0,
			o0 => Or227340_o0
		);
		Or227360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or227340_o0,
			i1 => And227200_o0,
			o0 => Or227360_o0
		);
		Or227380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or227360_o0,
			i1 => And227160_o0,
			o0 => Or227380_o0
		);
		And227400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12100_o0,
			i1 => i5,
			o0 => And227400_o0
		);
		And227420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23320_o0,
			i1 => i40,
			o0 => And227420_o0
		);
		And227440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227420_o0,
			i1 => And227400_o0,
			o0 => And227440_o0
		);
		And227460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227440_o0,
			i1 => Or227380_o0,
			o0 => And227460_o0
		);
		Or227480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227460_o0,
			i1 => And227000_o0,
			o0 => Or227480_o0
		);
		And227500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227480_o0,
			i1 => Not140_o0,
			o0 => And227500_o0
		);
		And227520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not540_o0,
			i1 => i3,
			o0 => And227520_o0
		);
		And227540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227520_o0,
			i1 => And226080_o0,
			o0 => And227540_o0
		);
		Or227560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227540_o0,
			i1 => And227500_o0,
			o0 => Or227560_o0
		);
		And227580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor226140_o0,
			i1 => Not3300_o0,
			o0 => And227580_o0
		);
		And227600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227580_o0,
			i1 => Nor23600_o0,
			o0 => And227600_o0
		);
		And227620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227600_o0,
			i1 => Or227560_o0,
			o0 => And227620_o0
		);
		And227640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220440_o0,
			i1 => Not12100_o0,
			o0 => And227640_o0
		);
		Or227660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227640_o0,
			i1 => And227620_o0,
			o0 => Or227660_o0
		);
		And227680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227660_o0,
			i1 => Not20520_o0,
			o0 => And227680_o0
		);
		Or227700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227680_o0,
			i1 => And226280_o0,
			o0 => Or227700_o0
		);
		Nor227720 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i31,
			i1 => i29,
			o0 => Nor227720_o0
		);
		And227740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216540_o0,
			i1 => i29,
			o0 => And227740_o0
		);
		Or227760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227740_o0,
			i1 => Nor227720_o0,
			o0 => Or227760_o0
		);
		And227780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227760_o0,
			i1 => Not80_o0,
			o0 => And227780_o0
		);
		Xor227800 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i17,
			o0 => Xor227800_o0
		);
		Not27820 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Xor227800_o0,
			o0 => Not27820_o0
		);
		And227840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not27820_o0,
			i1 => Nor26660_o0,
			o0 => And227840_o0
		);
		Or227860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => i16,
			o0 => Or227860_o0
		);
		Or227880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or227860_o0,
			i1 => And227840_o0,
			o0 => Or227880_o0
		);
		And227900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227880_o0,
			i1 => i14,
			o0 => And227900_o0
		);
		Or227920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227900_o0,
			i1 => And227780_o0,
			o0 => Or227920_o0
		);
		And227940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227920_o0,
			i1 => Not620_o0,
			o0 => And227940_o0
		);
		Or227960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226340_o0,
			i1 => i17,
			o0 => Or227960_o0
		);
		And227980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227960_o0,
			i1 => And28060_o0,
			o0 => And227980_o0
		);
		Or228000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227980_o0,
			i1 => And227940_o0,
			o0 => Or228000_o0
		);
		And228020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228000_o0,
			i1 => i13,
			o0 => And228020_o0
		);
		And228040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor216140_o0,
			i1 => i15,
			o0 => And228040_o0
		);
		Or228060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And212560_o0,
			i1 => And2240_o0,
			o0 => Or228060_o0
		);
		And228080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228060_o0,
			i1 => Not620_o0,
			o0 => And228080_o0
		);
		Or228100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228080_o0,
			i1 => And228040_o0,
			o0 => Or228100_o0
		);
		And228120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228100_o0,
			i1 => And210420_o0,
			o0 => And228120_o0
		);
		Xor228140 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i18,
			o0 => Xor228140_o0
		);
		Not28160 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Xor228140_o0,
			o0 => Not28160_o0
		);
		Or228180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i16,
			o0 => Or228180_o0
		);
		And228200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228180_o0,
			i1 => i15,
			o0 => And228200_o0
		);
		Or228220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228200_o0,
			i1 => And217280_o0,
			o0 => Or228220_o0
		);
		And228240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228220_o0,
			i1 => Not28160_o0,
			o0 => And228240_o0
		);
		And228260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1500_o0,
			i1 => i16,
			o0 => And228260_o0
		);
		And228280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228260_o0,
			i1 => i15,
			o0 => And228280_o0
		);
		Or228300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228280_o0,
			i1 => Xor2200_o0,
			o0 => Or228300_o0
		);
		And228320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228300_o0,
			i1 => i18,
			o0 => And228320_o0
		);
		And228340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215880_o0,
			i1 => Not620_o0,
			o0 => And228340_o0
		);
		Or228360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228340_o0,
			i1 => And22220_o0,
			o0 => Or228360_o0
		);
		And228380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228360_o0,
			i1 => Not1080_o0,
			o0 => And228380_o0
		);
		Or228400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228380_o0,
			i1 => And228320_o0,
			o0 => Or228400_o0
		);
		And228420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228400_o0,
			i1 => Not1040_o0,
			o0 => And228420_o0
		);
		Or228440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228420_o0,
			i1 => And228240_o0,
			o0 => Or228440_o0
		);
		Or228460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or228440_o0,
			i1 => And228120_o0,
			o0 => Or228460_o0
		);
		And228480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228460_o0,
			i1 => Not80_o0,
			o0 => And228480_o0
		);
		Or228500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228480_o0,
			i1 => And213180_o0,
			o0 => Or228500_o0
		);
		And228520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228500_o0,
			i1 => Not2080_o0,
			o0 => And228520_o0
		);
		Or228540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228520_o0,
			i1 => And228020_o0,
			o0 => Or228540_o0
		);
		And228560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228540_o0,
			i1 => i12,
			o0 => And228560_o0
		);
		And228580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i15,
			o0 => And228580_o0
		);
		And228600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228580_o0,
			i1 => And2240_o0,
			o0 => And228600_o0
		);
		Or228620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228600_o0,
			i1 => Not620_o0,
			o0 => Or228620_o0
		);
		And228640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228620_o0,
			i1 => And23520_o0,
			o0 => And228640_o0
		);
		And228660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223260_o0,
			i1 => And22300_o0,
			o0 => And228660_o0
		);
		And228680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => And22800_o0,
			o0 => And228680_o0
		);
		Or228700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228680_o0,
			i1 => And228660_o0,
			o0 => Or228700_o0
		);
		And228720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228700_o0,
			i1 => Not1080_o0,
			o0 => And228720_o0
		);
		And228740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => i17,
			o0 => And228740_o0
		);
		And228760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228740_o0,
			i1 => And226320_o0,
			o0 => And228760_o0
		);
		Or228780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228760_o0,
			i1 => And228720_o0,
			o0 => Or228780_o0
		);
		Or228800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or228780_o0,
			i1 => And228640_o0,
			o0 => Or228800_o0
		);
		And228820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228800_o0,
			i1 => Not1280_o0,
			o0 => And228820_o0
		);
		And228840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214100_o0,
			i1 => Not620_o0,
			o0 => And228840_o0
		);
		Or228860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228840_o0,
			i1 => And22800_o0,
			o0 => Or228860_o0
		);
		And228880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219620_o0,
			i1 => Not1080_o0,
			o0 => And228880_o0
		);
		And228900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228880_o0,
			i1 => Or228860_o0,
			o0 => And228900_o0
		);
		Or228920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228900_o0,
			i1 => i14,
			o0 => Or228920_o0
		);
		And228940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228920_o0,
			i1 => i13,
			o0 => And228940_o0
		);
		And228960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227020_o0,
			i1 => Not2080_o0,
			o0 => And228960_o0
		);
		And228980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => And2640_o0,
			o0 => And228980_o0
		);
		Or229000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228980_o0,
			i1 => And228960_o0,
			o0 => Or229000_o0
		);
		And229020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229000_o0,
			i1 => Not28160_o0,
			o0 => And229020_o0
		);
		And229040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219460_o0,
			i1 => Xor216140_o0,
			o0 => And229040_o0
		);
		And229060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => And2240_o0,
			o0 => And229060_o0
		);
		Or229080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229060_o0,
			i1 => And229040_o0,
			o0 => Or229080_o0
		);
		And229100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229080_o0,
			i1 => And223260_o0,
			o0 => And229100_o0
		);
		Or229120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229100_o0,
			i1 => And229020_o0,
			o0 => Or229120_o0
		);
		Or229140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or229120_o0,
			i1 => And228940_o0,
			o0 => Or229140_o0
		);
		Or229160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or229140_o0,
			i1 => And228820_o0,
			o0 => Or229160_o0
		);
		And229180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229160_o0,
			i1 => Not180_o0,
			o0 => And229180_o0
		);
		Or229200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229180_o0,
			i1 => And228560_o0,
			o0 => Or229200_o0
		);
		And229220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229200_o0,
			i1 => And26520_o0,
			o0 => And229220_o0
		);
		And229240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29680_o0,
			i1 => i22,
			o0 => And229240_o0
		);
		Or229260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229240_o0,
			i1 => And29820_o0,
			o0 => Or229260_o0
		);
		Nor229280 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			i1 => i19,
			o0 => Nor229280_o0
		);
		And229300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor229280_o0,
			i1 => i21,
			o0 => And229300_o0
		);
		And229320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => And21640_o0,
			o0 => And229320_o0
		);
		And229340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229320_o0,
			i1 => And23080_o0,
			o0 => And229340_o0
		);
		And229360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229340_o0,
			i1 => And229300_o0,
			o0 => And229360_o0
		);
		And229380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229360_o0,
			i1 => Or229260_o0,
			o0 => And229380_o0
		);
		Or229400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229380_o0,
			i1 => And211460_o0,
			o0 => Or229400_o0
		);
		And229420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i3,
			o0 => And229420_o0
		);
		And229440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229420_o0,
			i1 => Or229400_o0,
			o0 => And229440_o0
		);
		Or229460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229440_o0,
			i1 => And229220_o0,
			o0 => Or229460_o0
		);
		And229480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229460_o0,
			i1 => Not540_o0,
			o0 => And229480_o0
		);
		Nor229500 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor218020_o0,
			i1 => i22,
			o0 => Nor229500_o0
		);
		Or229520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor229500_o0,
			i1 => And221280_o0,
			o0 => Or229520_o0
		);
		And229540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229520_o0,
			i1 => And29560_o0,
			o0 => And229540_o0
		);
		Or229560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229540_o0,
			i1 => And218280_o0,
			o0 => Or229560_o0
		);
		And229580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => And22300_o0,
			o0 => And229580_o0
		);
		And229600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229580_o0,
			i1 => And23080_o0,
			o0 => And229600_o0
		);
		And229620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229600_o0,
			i1 => Or229560_o0,
			o0 => And229620_o0
		);
		Or229640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229620_o0,
			i1 => And211160_o0,
			o0 => Or229640_o0
		);
		And229660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229640_o0,
			i1 => Not1280_o0,
			o0 => And229660_o0
		);
		Or229680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229660_o0,
			i1 => And211360_o0,
			o0 => Or229680_o0
		);
		And229700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229680_o0,
			i1 => i3,
			o0 => And229700_o0
		);
		And229720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21520_o0,
			i1 => Not620_o0,
			o0 => And229720_o0
		);
		Or229740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229720_o0,
			i1 => And22800_o0,
			o0 => Or229740_o0
		);
		And229760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229740_o0,
			i1 => Not1080_o0,
			o0 => And229760_o0
		);
		Or229780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229760_o0,
			i1 => And22320_o0,
			o0 => Or229780_o0
		);
		And229800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229780_o0,
			i1 => i16,
			o0 => And229800_o0
		);
		And229820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226340_o0,
			i1 => i15,
			o0 => And229820_o0
		);
		Or229840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229820_o0,
			i1 => And229800_o0,
			o0 => Or229840_o0
		);
		And229860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224320_o0,
			i1 => Not180_o0,
			o0 => And229860_o0
		);
		And229880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229860_o0,
			i1 => Or229840_o0,
			o0 => And229880_o0
		);
		Or229900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229880_o0,
			i1 => And229700_o0,
			o0 => Or229900_o0
		);
		And229920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i5,
			o0 => And229920_o0
		);
		And229940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229920_o0,
			i1 => Or229900_o0,
			o0 => And229940_o0
		);
		Or229960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And229940_o0,
			i1 => And229480_o0,
			o0 => Or229960_o0
		);
		And229980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or229960_o0,
			i1 => Not160_o0,
			o0 => And229980_o0
		);
		And230000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217820_o0,
			i1 => Not540_o0,
			o0 => And230000_o0
		);
		Nor230020 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => i22,
			o0 => Nor230020_o0
		);
		And230040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor230020_o0,
			i1 => i5,
			o0 => And230040_o0
		);
		Or230060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230040_o0,
			i1 => And230000_o0,
			o0 => Or230060_o0
		);
		And230080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229600_o0,
			i1 => And210780_o0,
			o0 => And230080_o0
		);
		And230100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230080_o0,
			i1 => Or230060_o0,
			o0 => And230100_o0
		);
		Or230120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230100_o0,
			i1 => And211160_o0,
			o0 => Or230120_o0
		);
		And230140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230120_o0,
			i1 => Not1280_o0,
			o0 => And230140_o0
		);
		Or230160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230140_o0,
			i1 => And211360_o0,
			o0 => Or230160_o0
		);
		And230180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230160_o0,
			i1 => i3,
			o0 => And230180_o0
		);
		And230200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211460_o0,
			i1 => Not140_o0,
			o0 => And230200_o0
		);
		Or230220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230200_o0,
			i1 => And230180_o0,
			o0 => Or230220_o0
		);
		And230240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i4,
			o0 => And230240_o0
		);
		And230260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230240_o0,
			i1 => Or230220_o0,
			o0 => And230260_o0
		);
		Or230280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230260_o0,
			i1 => And229980_o0,
			o0 => Or230280_o0
		);
		And230300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230280_o0,
			i1 => Not120_o0,
			o0 => And230300_o0
		);
		And230320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222820_o0,
			i1 => i20,
			o0 => And230320_o0
		);
		And230340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230320_o0,
			i1 => And228740_o0,
			o0 => And230340_o0
		);
		And230360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => Not2080_o0,
			o0 => And230360_o0
		);
		And230380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22100_o0,
			i1 => Not140_o0,
			o0 => And230380_o0
		);
		And230400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230380_o0,
			i1 => And230360_o0,
			o0 => And230400_o0
		);
		And230420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230400_o0,
			i1 => And230340_o0,
			o0 => And230420_o0
		);
		Or230440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230420_o0,
			i1 => And211460_o0,
			o0 => Or230440_o0
		);
		And230460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor229280_o0,
			i1 => And21640_o0,
			o0 => And230460_o0
		);
		And230480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9800_o0,
			i1 => i21,
			o0 => And230480_o0
		);
		And230500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230480_o0,
			i1 => And221240_o0,
			o0 => And230500_o0
		);
		And230520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230500_o0,
			i1 => And230460_o0,
			o0 => And230520_o0
		);
		And230540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Nor21840_o0,
			o0 => And230540_o0
		);
		And230560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230540_o0,
			i1 => And24860_o0,
			o0 => And230560_o0
		);
		And230580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230560_o0,
			i1 => And230520_o0,
			o0 => And230580_o0
		);
		Or230600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230580_o0,
			i1 => Or230440_o0,
			o0 => Or230600_o0
		);
		And230620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i2,
			o0 => And230620_o0
		);
		And230640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230620_o0,
			i1 => Or230600_o0,
			o0 => And230640_o0
		);
		Or230660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230640_o0,
			i1 => And230300_o0,
			o0 => Or230660_o0
		);
		And230680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230660_o0,
			i1 => Not100_o0,
			o0 => And230680_o0
		);
		And230700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27500_o0,
			i1 => Not7440_o0,
			o0 => And230700_o0
		);
		And230720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21140_o0,
			i1 => Not160_o0,
			o0 => And230720_o0
		);
		And230740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230720_o0,
			i1 => And230700_o0,
			o0 => And230740_o0
		);
		And230760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => And22400_o0,
			o0 => And230760_o0
		);
		And230780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214860_o0,
			i1 => Nor21140_o0,
			o0 => And230780_o0
		);
		And230800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230780_o0,
			i1 => And230760_o0,
			o0 => And230800_o0
		);
		Or230820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230800_o0,
			i1 => And230740_o0,
			o0 => Or230820_o0
		);
		Or230840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or230820_o0,
			i1 => Or21020_o0,
			o0 => Or230840_o0
		);
		And230860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230840_o0,
			i1 => And223600_o0,
			o0 => And230860_o0
		);
		And230880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230860_o0,
			i1 => i1,
			o0 => And230880_o0
		);
		Or230900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And230880_o0,
			i1 => And230680_o0,
			o0 => Or230900_o0
		);
		And230920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230900_o0,
			i1 => Not60_o0,
			o0 => And230920_o0
		);
		Or230940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not140_o0,
			o0 => Or230940_o0
		);
		And230960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or230940_o0,
			i1 => Or22840_o0,
			o0 => And230960_o0
		);
		And230980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22800_o0,
			i1 => And21100_o0,
			o0 => And230980_o0
		);
		And231000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230980_o0,
			i1 => And24860_o0,
			o0 => And231000_o0
		);
		Or231020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231000_o0,
			i1 => And230960_o0,
			o0 => Or231020_o0
		);
		And231040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231020_o0,
			i1 => i16,
			o0 => And231040_o0
		);
		And231060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229820_o0,
			i1 => Nor21260_o0,
			o0 => And231060_o0
		);
		And231080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231060_o0,
			i1 => Not140_o0,
			o0 => And231080_o0
		);
		Or231100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231080_o0,
			i1 => And231040_o0,
			o0 => Or231100_o0
		);
		And231120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor27840_o0,
			i1 => And23520_o0,
			o0 => And231120_o0
		);
		And231140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231120_o0,
			i1 => And23180_o0,
			o0 => And231140_o0
		);
		And231160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231140_o0,
			i1 => Or231100_o0,
			o0 => And231160_o0
		);
		Or231180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231160_o0,
			i1 => And230920_o0,
			o0 => Or231180_o0
		);
		And231200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231180_o0,
			i1 => And23360_o0,
			o0 => And231200_o0
		);
		And231220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228740_o0,
			i1 => And23020_o0,
			o0 => And231220_o0
		);
		And231240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => And23080_o0,
			o0 => And231240_o0
		);
		And231260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210100_o0,
			i1 => And23020_o0,
			o0 => And231260_o0
		);
		Or231280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231260_o0,
			i1 => And231240_o0,
			o0 => Or231280_o0
		);
		Or231300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or231280_o0,
			i1 => And231220_o0,
			o0 => Or231300_o0
		);
		And231320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => And25600_o0,
			o0 => And231320_o0
		);
		And231340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231320_o0,
			i1 => And23340_o0,
			o0 => And231340_o0
		);
		And231360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231340_o0,
			i1 => And213280_o0,
			o0 => And231360_o0
		);
		And231380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231360_o0,
			i1 => Or231300_o0,
			o0 => And231380_o0
		);
		And231400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220920_o0,
			i1 => Not1500_o0,
			o0 => And231400_o0
		);
		And231420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231400_o0,
			i1 => And22300_o0,
			o0 => And231420_o0
		);
		And231440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29940_o0,
			i1 => i15,
			o0 => And231440_o0
		);
		Or231460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231440_o0,
			i1 => And231420_o0,
			o0 => Or231460_o0
		);
		And231480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231460_o0,
			i1 => Or210400_o0,
			o0 => And231480_o0
		);
		Or231500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i15,
			o0 => Or231500_o0
		);
		And231520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231500_o0,
			i1 => Not1500_o0,
			o0 => And231520_o0
		);
		And231540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29940_o0,
			i1 => Not620_o0,
			o0 => And231540_o0
		);
		Or231560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231540_o0,
			i1 => And231520_o0,
			o0 => Or231560_o0
		);
		And231580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231560_o0,
			i1 => Not540_o0,
			o0 => And231580_o0
		);
		And231600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214100_o0,
			i1 => And28460_o0,
			o0 => And231600_o0
		);
		Or231620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231600_o0,
			i1 => And231580_o0,
			o0 => Or231620_o0
		);
		And231640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231620_o0,
			i1 => i40,
			o0 => And231640_o0
		);
		Or231660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231640_o0,
			i1 => And231480_o0,
			o0 => Or231660_o0
		);
		And231680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231660_o0,
			i1 => i18,
			o0 => And231680_o0
		);
		Nand231700 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i37,
			o0 => Nand231700_o0
		);
		Or231720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand231700_o0,
			i1 => Not1040_o0,
			o0 => Or231720_o0
		);
		And231740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231720_o0,
			i1 => Not620_o0,
			o0 => And231740_o0
		);
		Or231760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231740_o0,
			i1 => And228580_o0,
			o0 => Or231760_o0
		);
		And231780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231760_o0,
			i1 => i19,
			o0 => And231780_o0
		);
		And231800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214120_o0,
			i1 => i15,
			o0 => And231800_o0
		);
		Or231820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231800_o0,
			i1 => And228840_o0,
			o0 => Or231820_o0
		);
		And231840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231820_o0,
			i1 => Not20760_o0,
			o0 => And231840_o0
		);
		Or231860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231840_o0,
			i1 => And226600_o0,
			o0 => Or231860_o0
		);
		Or231880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or231860_o0,
			i1 => And231780_o0,
			o0 => Or231880_o0
		);
		And231900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231880_o0,
			i1 => And2560_o0,
			o0 => And231900_o0
		);
		And231920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29200_o0,
			i1 => And21520_o0,
			o0 => And231920_o0
		);
		Or231940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231920_o0,
			i1 => And231900_o0,
			o0 => Or231940_o0
		);
		And231960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231940_o0,
			i1 => Not1080_o0,
			o0 => And231960_o0
		);
		Or231980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And231960_o0,
			i1 => And231680_o0,
			o0 => Or231980_o0
		);
		And232000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231980_o0,
			i1 => i12,
			o0 => And232000_o0
		);
		And232020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => Not180_o0,
			o0 => And232020_o0
		);
		Or232040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232020_o0,
			i1 => And232000_o0,
			o0 => Or232040_o0
		);
		And232060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232040_o0,
			i1 => Not1280_o0,
			o0 => And232060_o0
		);
		Nand232080 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => Not1500_o0,
			o0 => Nand232080_o0
		);
		And232100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand232080_o0,
			i1 => Not1080_o0,
			o0 => And232100_o0
		);
		Or232120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232100_o0,
			i1 => And215060_o0,
			o0 => Or232120_o0
		);
		And232140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222800_o0,
			i1 => And22300_o0,
			o0 => And232140_o0
		);
		And232160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And232140_o0,
			i1 => Or232120_o0,
			o0 => And232160_o0
		);
		And232180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => Not620_o0,
			o0 => And232180_o0
		);
		And232200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And232180_o0,
			i1 => And222800_o0,
			o0 => And232200_o0
		);
		Nor232220 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i5,
			o0 => Nor232220_o0
		);
		And232240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213520_o0,
			i1 => i5,
			o0 => And232240_o0
		);
		Or232260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232240_o0,
			i1 => Nor232220_o0,
			o0 => Or232260_o0
		);
		Or232280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or232260_o0,
			i1 => And232200_o0,
			o0 => Or232280_o0
		);
		Or232300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or232280_o0,
			i1 => And232160_o0,
			o0 => Or232300_o0
		);
		And232320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232300_o0,
			i1 => And28480_o0,
			o0 => And232320_o0
		);
		Or232340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232320_o0,
			i1 => And232060_o0,
			o0 => Or232340_o0
		);
		And232360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232340_o0,
			i1 => Not80_o0,
			o0 => And232360_o0
		);
		And232380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219480_o0,
			i1 => i5,
			o0 => And232380_o0
		);
		And232400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226340_o0,
			i1 => Nor21980_o0,
			o0 => And232400_o0
		);
		And232420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => Not540_o0,
			o0 => And232420_o0
		);
		And232440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And232420_o0,
			i1 => And215080_o0,
			o0 => And232440_o0
		);
		Or232460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232440_o0,
			i1 => And232400_o0,
			o0 => Or232460_o0
		);
		Or232480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or232460_o0,
			i1 => And232380_o0,
			o0 => Or232480_o0
		);
		And232500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232480_o0,
			i1 => Not180_o0,
			o0 => And232500_o0
		);
		And232520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213520_o0,
			i1 => Not540_o0,
			o0 => And232520_o0
		);
		Or232540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232520_o0,
			i1 => And232500_o0,
			o0 => Or232540_o0
		);
		And232560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232540_o0,
			i1 => And24040_o0,
			o0 => And232560_o0
		);
		Or232580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232560_o0,
			i1 => And232360_o0,
			o0 => Or232580_o0
		);
		And232600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232580_o0,
			i1 => Not2080_o0,
			o0 => And232600_o0
		);
		Not32620 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => i29,
			o0 => Not32620_o0
		);
		And232640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not32620_o0,
			i1 => i12,
			o0 => And232640_o0
		);
		And232660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor216140_o0,
			i1 => Not1040_o0,
			o0 => And232660_o0
		);
		Or232680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232660_o0,
			i1 => And228740_o0,
			o0 => Or232680_o0
		);
		And232700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232680_o0,
			i1 => And24880_o0,
			o0 => And232700_o0
		);
		Or232720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232700_o0,
			i1 => And232640_o0,
			o0 => Or232720_o0
		);
		And232740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232720_o0,
			i1 => Not620_o0,
			o0 => And232740_o0
		);
		And232760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223960_o0,
			i1 => i16,
			o0 => And232760_o0
		);
		Or232780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232760_o0,
			i1 => And212900_o0,
			o0 => Or232780_o0
		);
		Or232800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or232780_o0,
			i1 => i12,
			o0 => Or232800_o0
		);
		And232820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232800_o0,
			i1 => i15,
			o0 => And232820_o0
		);
		Or232840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232820_o0,
			i1 => And232740_o0,
			o0 => Or232840_o0
		);
		And232860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232840_o0,
			i1 => Not80_o0,
			o0 => And232860_o0
		);
		And232880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => And21100_o0,
			o0 => And232880_o0
		);
		Or232900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And26580_o0,
			i1 => i15,
			o0 => Or232900_o0
		);
		Or232920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or232900_o0,
			i1 => And232880_o0,
			o0 => Or232920_o0
		);
		And232940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232920_o0,
			i1 => Not1040_o0,
			o0 => And232940_o0
		);
		Or232960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232940_o0,
			i1 => And23060_o0,
			o0 => Or232960_o0
		);
		And232980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or232960_o0,
			i1 => i12,
			o0 => And232980_o0
		);
		And233000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not180_o0,
			o0 => And233000_o0
		);
		Or233020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233000_o0,
			i1 => And232980_o0,
			o0 => Or233020_o0
		);
		And233040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233020_o0,
			i1 => i14,
			o0 => And233040_o0
		);
		Or233060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233040_o0,
			i1 => And232860_o0,
			o0 => Or233060_o0
		);
		And233080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233060_o0,
			i1 => Not540_o0,
			o0 => And233080_o0
		);
		And233100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => And2640_o0,
			o0 => And233100_o0
		);
		Or233120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227280_o0,
			i1 => And227220_o0,
			o0 => Or233120_o0
		);
		Or233140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or233120_o0,
			i1 => And233100_o0,
			o0 => Or233140_o0
		);
		And233160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211020_o0,
			i1 => i14,
			o0 => And233160_o0
		);
		And233180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233160_o0,
			i1 => Or233140_o0,
			o0 => And233180_o0
		);
		Or233200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233180_o0,
			i1 => And233080_o0,
			o0 => Or233200_o0
		);
		And233220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233200_o0,
			i1 => i40,
			o0 => And233220_o0
		);
		And233240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226000_o0,
			i1 => And24280_o0,
			o0 => And233240_o0
		);
		Or233260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233240_o0,
			i1 => And233220_o0,
			o0 => Or233260_o0
		);
		And233280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233260_o0,
			i1 => i13,
			o0 => And233280_o0
		);
		Nor233300 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i5,
			o0 => Nor233300_o0
		);
		Or233320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor233300_o0,
			i1 => And233280_o0,
			o0 => Or233320_o0
		);
		Or233340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or233320_o0,
			i1 => And232600_o0,
			o0 => Or233340_o0
		);
		And233360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233340_o0,
			i1 => Not160_o0,
			o0 => And233360_o0
		);
		And233380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29940_o0,
			i1 => And23080_o0,
			o0 => And233380_o0
		);
		And233400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And21520_o0,
			o0 => And233400_o0
		);
		Or233420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233400_o0,
			i1 => And233380_o0,
			o0 => Or233420_o0
		);
		And233440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233420_o0,
			i1 => i18,
			o0 => And233440_o0
		);
		Or233460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233440_o0,
			i1 => And231260_o0,
			o0 => Or233460_o0
		);
		And233480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233460_o0,
			i1 => i15,
			o0 => And233480_o0
		);
		And233500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22300_o0,
			i1 => Not1500_o0,
			o0 => And233500_o0
		);
		And233520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233500_o0,
			i1 => And23080_o0,
			o0 => And233520_o0
		);
		And233540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233520_o0,
			i1 => Or221040_o0,
			o0 => And233540_o0
		);
		Or233560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233540_o0,
			i1 => And233480_o0,
			o0 => Or233560_o0
		);
		And233580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230240_o0,
			i1 => Not1280_o0,
			o0 => And233580_o0
		);
		And233600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233580_o0,
			i1 => Or233560_o0,
			o0 => And233600_o0
		);
		Or233620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233600_o0,
			i1 => And233360_o0,
			o0 => Or233620_o0
		);
		And233640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233620_o0,
			i1 => Not140_o0,
			o0 => And233640_o0
		);
		And233660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225320_o0,
			i1 => Not180_o0,
			o0 => And233660_o0
		);
		And233680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210660_o0,
			i1 => i22,
			o0 => And233680_o0
		);
		Or233700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233680_o0,
			i1 => And210740_o0,
			o0 => Or233700_o0
		);
		And233720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233700_o0,
			i1 => i27,
			o0 => And233720_o0
		);
		And233740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233720_o0,
			i1 => And29560_o0,
			o0 => And233740_o0
		);
		And233760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9700_o0,
			i1 => i22,
			o0 => And233760_o0
		);
		Or233780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor230020_o0,
			i1 => And233760_o0,
			o0 => Or233780_o0
		);
		And233800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233780_o0,
			i1 => And29560_o0,
			o0 => And233800_o0
		);
		Or233820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233800_o0,
			i1 => And210540_o0,
			o0 => Or233820_o0
		);
		Or233840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or233820_o0,
			i1 => And233740_o0,
			o0 => Or233840_o0
		);
		Or233860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or233840_o0,
			i1 => Not1080_o0,
			o0 => Or233860_o0
		);
		And233880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233860_o0,
			i1 => And211240_o0,
			o0 => And233880_o0
		);
		Or233900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233880_o0,
			i1 => And233660_o0,
			o0 => Or233900_o0
		);
		And233920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233900_o0,
			i1 => Not540_o0,
			o0 => And233920_o0
		);
		And233940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221200_o0,
			i1 => And233760_o0,
			o0 => And233940_o0
		);
		And233960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221240_o0,
			i1 => Not9800_o0,
			o0 => And233960_o0
		);
		Or233980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233960_o0,
			i1 => And233940_o0,
			o0 => Or233980_o0
		);
		And234000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or233980_o0,
			i1 => And29560_o0,
			o0 => And234000_o0
		);
		Or234020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234000_o0,
			i1 => And230320_o0,
			o0 => Or234020_o0
		);
		And234040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => i18,
			o0 => And234040_o0
		);
		And234060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234040_o0,
			i1 => And211020_o0,
			o0 => And234060_o0
		);
		And234080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234060_o0,
			i1 => Or234020_o0,
			o0 => And234080_o0
		);
		Or234100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234080_o0,
			i1 => And233920_o0,
			o0 => Or234100_o0
		);
		And234120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or234100_o0,
			i1 => Not160_o0,
			o0 => And234120_o0
		);
		Nor234140 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			i1 => i5,
			o0 => Nor234140_o0
		);
		And234160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor230020_o0,
			i1 => i21,
			o0 => And234160_o0
		);
		And234180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234160_o0,
			i1 => Nor234140_o0,
			o0 => And234180_o0
		);
		And234200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210580_o0,
			i1 => And233760_o0,
			o0 => And234200_o0
		);
		Or234220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234200_o0,
			i1 => And210540_o0,
			o0 => Or234220_o0
		);
		Or234240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or234220_o0,
			i1 => And234180_o0,
			o0 => Or234240_o0
		);
		And234260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i12,
			o0 => And234260_o0
		);
		And234280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234260_o0,
			i1 => Nor211040_o0,
			o0 => And234280_o0
		);
		And234300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234280_o0,
			i1 => And222240_o0,
			o0 => And234300_o0
		);
		And234320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234300_o0,
			i1 => Or234240_o0,
			o0 => And234320_o0
		);
		Or234340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234320_o0,
			i1 => And234120_o0,
			o0 => Or234340_o0
		);
		And234360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or234340_o0,
			i1 => Not1500_o0,
			o0 => And234360_o0
		);
		And234380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => Not160_o0,
			o0 => And234380_o0
		);
		And234400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor232220_o0,
			i1 => And225320_o0,
			o0 => And234400_o0
		);
		And234420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234400_o0,
			i1 => And234380_o0,
			o0 => And234420_o0
		);
		Or234440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234420_o0,
			i1 => And234360_o0,
			o0 => Or234440_o0
		);
		And234460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229420_o0,
			i1 => And21940_o0,
			o0 => And234460_o0
		);
		And234480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234460_o0,
			i1 => Or234440_o0,
			o0 => And234480_o0
		);
		Or234500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234480_o0,
			i1 => And233640_o0,
			o0 => Or234500_o0
		);
		And234520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or234500_o0,
			i1 => Not120_o0,
			o0 => And234520_o0
		);
		And234540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			i1 => i21,
			o0 => And234540_o0
		);
		And234560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221240_o0,
			i1 => Not9700_o0,
			o0 => And234560_o0
		);
		And234580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234560_o0,
			i1 => And234540_o0,
			o0 => And234580_o0
		);
		And234600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234580_o0,
			i1 => And230460_o0,
			o0 => And234600_o0
		);
		And234620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214660_o0,
			i1 => And23080_o0,
			o0 => And234620_o0
		);
		And234640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219060_o0,
			i1 => Nor21260_o0,
			o0 => And234640_o0
		);
		And234660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234640_o0,
			i1 => And234620_o0,
			o0 => And234660_o0
		);
		And234680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234660_o0,
			i1 => And234600_o0,
			o0 => And234680_o0
		);
		Or234700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234680_o0,
			i1 => And234520_o0,
			o0 => Or234700_o0
		);
		And234720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or234700_o0,
			i1 => Not60_o0,
			o0 => And234720_o0
		);
		And234740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214620_o0,
			i1 => Nor21140_o0,
			o0 => And234740_o0
		);
		And234760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234740_o0,
			i1 => And222800_o0,
			o0 => And234760_o0
		);
		And234780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => Not2080_o0,
			o0 => And234780_o0
		);
		And234800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234780_o0,
			i1 => And21960_o0,
			o0 => And234800_o0
		);
		And234820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234800_o0,
			i1 => And234760_o0,
			o0 => And234820_o0
		);
		Or234840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234820_o0,
			i1 => And234720_o0,
			o0 => Or234840_o0
		);
		Nor234860 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i1,
			o0 => Nor234860_o0
		);
		And234880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor234860_o0,
			i1 => Or234840_o0,
			o0 => And234880_o0
		);
		Or234900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234880_o0,
			i1 => i36,
			o0 => Or234900_o0
		);
		Or234920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or234900_o0,
			i1 => i10,
			o0 => Or234920_o0
		);
		Or234940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or234920_o0,
			i1 => i9,
			o0 => Or234940_o0
		);
		And234960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or234940_o0,
			i1 => Not24960_o0,
			o0 => And234960_o0
		);
		Or234980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => i9,
			o0 => Or234980_o0
		);
		And235000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or234980_o0,
			i1 => i11,
			o0 => And235000_o0
		);
		Or235020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235000_o0,
			i1 => And234960_o0,
			o0 => Or235020_o0
		);
		And235040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235020_o0,
			i1 => Not12100_o0,
			o0 => And235040_o0
		);
		And235060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220540_o0,
			i1 => Not20520_o0,
			o0 => And235060_o0
		);
		And235080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235060_o0,
			i1 => And23640_o0,
			o0 => And235080_o0
		);
		Or235100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235080_o0,
			i1 => And235040_o0,
			o0 => Or235100_o0
		);
		Nand235120 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			i1 => i20,
			o0 => Nand235120_o0
		);
		Or235140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand235120_o0,
			i1 => Not32620_o0,
			o0 => Or235140_o0
		);
		And235160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235140_o0,
			i1 => And23900_o0,
			o0 => And235160_o0
		);
		And235180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => i18,
			o0 => And235180_o0
		);
		And235200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => Not1080_o0,
			o0 => And235200_o0
		);
		Or235220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235200_o0,
			i1 => And235180_o0,
			o0 => Or235220_o0
		);
		And235240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21300_o0,
			i1 => Not1040_o0,
			o0 => And235240_o0
		);
		And235260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235240_o0,
			i1 => Or235220_o0,
			o0 => And235260_o0
		);
		Or235280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235260_o0,
			i1 => And235160_o0,
			o0 => Or235280_o0
		);
		And235300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235280_o0,
			i1 => i12,
			o0 => And235300_o0
		);
		And235320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28060_o0,
			i1 => And23020_o0,
			o0 => And235320_o0
		);
		Or235340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235320_o0,
			i1 => And235300_o0,
			o0 => Or235340_o0
		);
		And235360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235340_o0,
			i1 => And213300_o0,
			o0 => And235360_o0
		);
		And235380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210400_o0,
			i1 => Not120_o0,
			o0 => And235380_o0
		);
		And235400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not540_o0,
			i1 => i2,
			o0 => And235400_o0
		);
		And235420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235400_o0,
			i1 => And221240_o0,
			o0 => And235420_o0
		);
		Or235440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235420_o0,
			i1 => And235380_o0,
			o0 => Or235440_o0
		);
		And235460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235440_o0,
			i1 => Nand210560_o0,
			o0 => And235460_o0
		);
		And235480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			i1 => Not120_o0,
			o0 => And235480_o0
		);
		And235500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235480_o0,
			i1 => i23,
			o0 => And235500_o0
		);
		And235520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235500_o0,
			i1 => Or210400_o0,
			o0 => And235520_o0
		);
		Or235540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235520_o0,
			i1 => And235460_o0,
			o0 => Or235540_o0
		);
		And235560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235540_o0,
			i1 => Not9540_o0,
			o0 => And235560_o0
		);
		And235580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			i1 => Not120_o0,
			o0 => And235580_o0
		);
		And235600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235580_o0,
			i1 => Or210400_o0,
			o0 => And235600_o0
		);
		Or235620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235600_o0,
			i1 => And235560_o0,
			o0 => Or235620_o0
		);
		And235640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235620_o0,
			i1 => i21,
			o0 => And235640_o0
		);
		And235660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235580_o0,
			i1 => Not10520_o0,
			o0 => And235660_o0
		);
		And235680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235660_o0,
			i1 => Or210400_o0,
			o0 => And235680_o0
		);
		Or235700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235680_o0,
			i1 => And235640_o0,
			o0 => Or235700_o0
		);
		And235720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235700_o0,
			i1 => i18,
			o0 => And235720_o0
		);
		And235740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => Not120_o0,
			o0 => And235740_o0
		);
		And235760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235740_o0,
			i1 => Not1080_o0,
			o0 => And235760_o0
		);
		Or235780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235760_o0,
			i1 => And235720_o0,
			o0 => Or235780_o0
		);
		And235800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235780_o0,
			i1 => Not1500_o0,
			o0 => And235800_o0
		);
		Nor235820 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i2,
			o0 => Nor235820_o0
		);
		And235840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor235820_o0,
			i1 => And224600_o0,
			o0 => And235840_o0
		);
		Or235860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235840_o0,
			i1 => And235800_o0,
			o0 => Or235860_o0
		);
		And235880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235860_o0,
			i1 => i17,
			o0 => And235880_o0
		);
		And235900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor235820_o0,
			i1 => And28040_o0,
			o0 => And235900_o0
		);
		And235920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And235900_o0,
			i1 => Or21720_o0,
			o0 => And235920_o0
		);
		Or235940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And235920_o0,
			i1 => And235880_o0,
			o0 => Or235940_o0
		);
		And235960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235940_o0,
			i1 => Not620_o0,
			o0 => And235960_o0
		);
		Or235980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not1040_o0,
			o0 => Or235980_o0
		);
		And236000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i5,
			o0 => And236000_o0
		);
		And236020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236000_o0,
			i1 => Or235980_o0,
			o0 => And236020_o0
		);
		And236040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not540_o0,
			o0 => And236040_o0
		);
		And236060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236040_o0,
			i1 => And222120_o0,
			o0 => And236060_o0
		);
		Or236080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236060_o0,
			i1 => And236020_o0,
			o0 => Or236080_o0
		);
		And236100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236080_o0,
			i1 => i18,
			o0 => And236100_o0
		);
		And236120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => Not1080_o0,
			o0 => And236120_o0
		);
		And236140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236120_o0,
			i1 => Not27820_o0,
			o0 => And236140_o0
		);
		Or236160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236140_o0,
			i1 => And236100_o0,
			o0 => Or236160_o0
		);
		And236180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not120_o0,
			o0 => And236180_o0
		);
		And236200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236180_o0,
			i1 => Or236160_o0,
			o0 => And236200_o0
		);
		Or236220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236200_o0,
			i1 => And235960_o0,
			o0 => Or236220_o0
		);
		And236240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236220_o0,
			i1 => i12,
			o0 => And236240_o0
		);
		And236260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And232020_o0,
			i1 => Not120_o0,
			o0 => And236260_o0
		);
		Or236280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236260_o0,
			i1 => And236240_o0,
			o0 => Or236280_o0
		);
		And236300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236280_o0,
			i1 => Not1280_o0,
			o0 => And236300_o0
		);
		And236320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And232320_o0,
			i1 => Not120_o0,
			o0 => And236320_o0
		);
		Or236340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236320_o0,
			i1 => And236300_o0,
			o0 => Or236340_o0
		);
		And236360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236340_o0,
			i1 => Not2080_o0,
			o0 => And236360_o0
		);
		Nor236380 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor26980_o0,
			i1 => Not540_o0,
			o0 => Nor236380_o0
		);
		Nor236400 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i5,
			o0 => Nor236400_o0
		);
		And236420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor236400_o0,
			i1 => And24940_o0,
			o0 => And236420_o0
		);
		Or236440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236420_o0,
			i1 => Nor236380_o0,
			o0 => Or236440_o0
		);
		And236460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236440_o0,
			i1 => And21300_o0,
			o0 => And236460_o0
		);
		Or236480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236460_o0,
			i1 => And216060_o0,
			o0 => Or236480_o0
		);
		And236500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236480_o0,
			i1 => Not1500_o0,
			o0 => And236500_o0
		);
		And236520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210100_o0,
			i1 => i15,
			o0 => And236520_o0
		);
		Xor236540 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => Not620_o0,
			o0 => Xor236540_o0
		);
		Or236560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Xor236540_o0,
			i1 => And236520_o0,
			o0 => Or236560_o0
		);
		And236580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236560_o0,
			i1 => i16,
			o0 => And236580_o0
		);
		And236600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223960_o0,
			i1 => And21300_o0,
			o0 => And236600_o0
		);
		Or236620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236600_o0,
			i1 => And236580_o0,
			o0 => Or236620_o0
		);
		And236640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236620_o0,
			i1 => And2560_o0,
			o0 => And236640_o0
		);
		And236660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224160_o0,
			i1 => And28460_o0,
			o0 => And236660_o0
		);
		And236680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => i19,
			o0 => And236680_o0
		);
		And236700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236680_o0,
			i1 => And22400_o0,
			o0 => And236700_o0
		);
		And236720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236700_o0,
			i1 => Or210400_o0,
			o0 => And236720_o0
		);
		Or236740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236720_o0,
			i1 => And236660_o0,
			o0 => Or236740_o0
		);
		Or236760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or236740_o0,
			i1 => And236640_o0,
			o0 => Or236760_o0
		);
		Or236780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or236760_o0,
			i1 => And236500_o0,
			o0 => Or236780_o0
		);
		And236800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or236780_o0,
			i1 => Not180_o0,
			o0 => And236800_o0
		);
		And236820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i29,
			i1 => i23,
			o0 => And236820_o0
		);
		Nor236840 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			i1 => i15,
			o0 => Nor236840_o0
		);
		And236860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor236840_o0,
			i1 => And216540_o0,
			o0 => And236860_o0
		);
		And236880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236860_o0,
			i1 => And236820_o0,
			o0 => And236880_o0
		);
		Or236900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236880_o0,
			i1 => i15,
			o0 => Or236900_o0
		);
		And236920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222800_o0,
			i1 => i40,
			o0 => And236920_o0
		);
		And236940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236920_o0,
			i1 => Or236900_o0,
			o0 => And236940_o0
		);
		Or236960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And236940_o0,
			i1 => And236800_o0,
			o0 => Or236960_o0
		);
		And236980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => Not120_o0,
			o0 => And236980_o0
		);
		And237000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236980_o0,
			i1 => Or236960_o0,
			o0 => And237000_o0
		);
		Or237020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237000_o0,
			i1 => And236360_o0,
			o0 => Or237020_o0
		);
		And237040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237020_o0,
			i1 => Not140_o0,
			o0 => And237040_o0
		);
		And237060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233760_o0,
			i1 => i18,
			o0 => And237060_o0
		);
		And237080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29720_o0,
			i1 => And29560_o0,
			o0 => And237080_o0
		);
		And237100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237080_o0,
			i1 => And237060_o0,
			o0 => And237100_o0
		);
		Or237120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237100_o0,
			i1 => Not1080_o0,
			o0 => Or237120_o0
		);
		And237140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237120_o0,
			i1 => And211240_o0,
			o0 => And237140_o0
		);
		Or237160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237140_o0,
			i1 => And233660_o0,
			o0 => Or237160_o0
		);
		And237180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237160_o0,
			i1 => Not1500_o0,
			o0 => And237180_o0
		);
		And237200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => i15,
			o0 => And237200_o0
		);
		And237220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237200_o0,
			i1 => And23020_o0,
			o0 => And237220_o0
		);
		Or237240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237220_o0,
			i1 => And237180_o0,
			o0 => Or237240_o0
		);
		And237260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236040_o0,
			i1 => Not1280_o0,
			o0 => And237260_o0
		);
		And237280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237260_o0,
			i1 => And26040_o0,
			o0 => And237280_o0
		);
		And237300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237280_o0,
			i1 => Or237240_o0,
			o0 => And237300_o0
		);
		Or237320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237300_o0,
			i1 => And237040_o0,
			o0 => Or237320_o0
		);
		And237340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237320_o0,
			i1 => Not60_o0,
			o0 => And237340_o0
		);
		And237360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229820_o0,
			i1 => Not140_o0,
			o0 => And237360_o0
		);
		Or237380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237360_o0,
			i1 => And218640_o0,
			o0 => Or237380_o0
		);
		And237400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237380_o0,
			i1 => And23020_o0,
			o0 => And237400_o0
		);
		Or237420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237400_o0,
			i1 => And218760_o0,
			o0 => Or237420_o0
		);
		And237440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not120_o0,
			i1 => i0,
			o0 => And237440_o0
		);
		And237460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237440_o0,
			i1 => Not540_o0,
			o0 => And237460_o0
		);
		And237480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237460_o0,
			i1 => Or237420_o0,
			o0 => And237480_o0
		);
		Or237500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237480_o0,
			i1 => And237340_o0,
			o0 => Or237500_o0
		);
		And237520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237500_o0,
			i1 => Not100_o0,
			o0 => And237520_o0
		);
		And237540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224460_o0,
			i1 => And21300_o0,
			o0 => And237540_o0
		);
		And237560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237540_o0,
			i1 => Nor232220_o0,
			o0 => And237560_o0
		);
		Nor237580 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i3,
			i1 => i0,
			o0 => Nor237580_o0
		);
		And237600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor237580_o0,
			i1 => i13,
			o0 => And237600_o0
		);
		And237620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237600_o0,
			i1 => And21240_o0,
			o0 => And237620_o0
		);
		And237640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237620_o0,
			i1 => And237560_o0,
			o0 => And237640_o0
		);
		Or237660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237640_o0,
			i1 => And237520_o0,
			o0 => Or237660_o0
		);
		And237680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237660_o0,
			i1 => Not160_o0,
			o0 => And237680_o0
		);
		Xor237700 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i3,
			o0 => Xor237700_o0
		);
		And237720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215240_o0,
			i1 => And211240_o0,
			o0 => And237720_o0
		);
		Or237740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237720_o0,
			i1 => And211160_o0,
			o0 => Or237740_o0
		);
		And237760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237740_o0,
			i1 => Not1280_o0,
			o0 => And237760_o0
		);
		Or237780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237760_o0,
			i1 => And211360_o0,
			o0 => Or237780_o0
		);
		And237800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237780_o0,
			i1 => Not120_o0,
			o0 => And237800_o0
		);
		Or237820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237800_o0,
			i1 => And211540_o0,
			o0 => Or237820_o0
		);
		And237840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237820_o0,
			i1 => Not100_o0,
			o0 => And237840_o0
		);
		And237860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Or21020_o0,
			o0 => And237860_o0
		);
		And237880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237860_o0,
			i1 => i1,
			o0 => And237880_o0
		);
		Or237900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And237880_o0,
			i1 => And237840_o0,
			o0 => Or237900_o0
		);
		And237920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or237900_o0,
			i1 => Xor237700_o0,
			o0 => And237920_o0
		);
		And237940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not140_o0,
			o0 => And237940_o0
		);
		And237960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237940_o0,
			i1 => Not120_o0,
			o0 => And237960_o0
		);
		And237980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i3,
			i1 => i2,
			o0 => And237980_o0
		);
		And238000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237980_o0,
			i1 => Not1040_o0,
			o0 => And238000_o0
		);
		Or238020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238000_o0,
			i1 => And237960_o0,
			o0 => Or238020_o0
		);
		And238040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238020_o0,
			i1 => Not1080_o0,
			o0 => And238040_o0
		);
		And238060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228740_o0,
			i1 => Nor21140_o0,
			o0 => And238060_o0
		);
		Or238080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238060_o0,
			i1 => And238040_o0,
			o0 => Or238080_o0
		);
		And238100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238080_o0,
			i1 => And23020_o0,
			o0 => And238100_o0
		);
		Nor238120 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i13,
			o0 => Nor238120_o0
		);
		And238140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor238120_o0,
			i1 => And2240_o0,
			o0 => And238140_o0
		);
		And238160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238140_o0,
			i1 => And24160_o0,
			o0 => And238160_o0
		);
		Or238180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238160_o0,
			i1 => And238100_o0,
			o0 => Or238180_o0
		);
		And238200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238180_o0,
			i1 => i15,
			o0 => And238200_o0
		);
		And238220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221240_o0,
			i1 => i3,
			o0 => And238220_o0
		);
		And238240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29720_o0,
			i1 => Not140_o0,
			o0 => And238240_o0
		);
		Or238260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238240_o0,
			i1 => And238220_o0,
			o0 => Or238260_o0
		);
		And238280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238260_o0,
			i1 => Nand210560_o0,
			o0 => And238280_o0
		);
		And238300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229240_o0,
			i1 => Not140_o0,
			o0 => And238300_o0
		);
		Or238320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238300_o0,
			i1 => And238280_o0,
			o0 => Or238320_o0
		);
		And238340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9540_o0,
			i1 => i18,
			o0 => And238340_o0
		);
		And238360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238340_o0,
			i1 => i21,
			o0 => And238360_o0
		);
		And238380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238360_o0,
			i1 => Or238320_o0,
			o0 => And238380_o0
		);
		Nor238400 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i3,
			o0 => Nor238400_o0
		);
		Or238420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor238400_o0,
			i1 => And238380_o0,
			o0 => Or238420_o0
		);
		And238440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => Not120_o0,
			o0 => And238440_o0
		);
		And238460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => And21520_o0,
			o0 => And238460_o0
		);
		And238480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238460_o0,
			i1 => And238440_o0,
			o0 => And238480_o0
		);
		And238500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238480_o0,
			i1 => Or238420_o0,
			o0 => And238500_o0
		);
		Or238520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238500_o0,
			i1 => And238200_o0,
			o0 => Or238520_o0
		);
		And238540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238520_o0,
			i1 => Not1280_o0,
			o0 => And238540_o0
		);
		And238560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237980_o0,
			i1 => And211360_o0,
			o0 => And238560_o0
		);
		Or238580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238560_o0,
			i1 => And238540_o0,
			o0 => Or238580_o0
		);
		And238600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238580_o0,
			i1 => Not100_o0,
			o0 => And238600_o0
		);
		And238620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i2,
			i1 => i1,
			o0 => And238620_o0
		);
		And238640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238620_o0,
			i1 => i3,
			o0 => And238640_o0
		);
		And238660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238640_o0,
			i1 => And237860_o0,
			o0 => And238660_o0
		);
		Or238680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238660_o0,
			i1 => And238600_o0,
			o0 => Or238680_o0
		);
		And238700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238680_o0,
			i1 => i4,
			o0 => And238700_o0
		);
		And238720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26040_o0,
			i1 => i4,
			o0 => And238720_o0
		);
		And238740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22600_o0,
			i1 => i2,
			o0 => And238740_o0
		);
		Or238760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238740_o0,
			i1 => And238720_o0,
			o0 => Or238760_o0
		);
		And238780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230700_o0,
			i1 => Not100_o0,
			o0 => And238780_o0
		);
		Or238800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238780_o0,
			i1 => Or21020_o0,
			o0 => Or238800_o0
		);
		And238820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238800_o0,
			i1 => And23020_o0,
			o0 => And238820_o0
		);
		And238840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230360_o0,
			i1 => And217160_o0,
			o0 => And238840_o0
		);
		And238860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238840_o0,
			i1 => And230340_o0,
			o0 => And238860_o0
		);
		Or238880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238860_o0,
			i1 => And238820_o0,
			o0 => Or238880_o0
		);
		And238900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238880_o0,
			i1 => Or238760_o0,
			o0 => And238900_o0
		);
		Or238920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i16,
			o0 => Or238920_o0
		);
		And238940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or238920_o0,
			i1 => And27500_o0,
			o0 => And238940_o0
		);
		Or238960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And238940_o0,
			i1 => And2660_o0,
			o0 => Or238960_o0
		);
		And238980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Nor22600_o0,
			o0 => And238980_o0
		);
		And239000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238980_o0,
			i1 => And224460_o0,
			o0 => And239000_o0
		);
		And239020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239000_o0,
			i1 => Or238960_o0,
			o0 => And239020_o0
		);
		Or239040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239020_o0,
			i1 => And238900_o0,
			o0 => Or239040_o0
		);
		Or239060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239040_o0,
			i1 => And238700_o0,
			o0 => Or239060_o0
		);
		Or239080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239060_o0,
			i1 => And237920_o0,
			o0 => Or239080_o0
		);
		And239100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239080_o0,
			i1 => Not60_o0,
			o0 => And239100_o0
		);
		And239120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And22860_o0,
			o0 => And239120_o0
		);
		And239140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239120_o0,
			i1 => And211740_o0,
			o0 => And239140_o0
		);
		Or239160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239140_o0,
			i1 => And239100_o0,
			o0 => Or239160_o0
		);
		Or239180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239160_o0,
			i1 => And237680_o0,
			o0 => Or239180_o0
		);
		And239200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239180_o0,
			i1 => Not80_o0,
			o0 => And239200_o0
		);
		Xor239220 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i17,
			o0 => Xor239220_o0
		);
		And239240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225220_o0,
			i1 => Nor26660_o0,
			o0 => And239240_o0
		);
		And239260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239240_o0,
			i1 => Xor239220_o0,
			o0 => And239260_o0
		);
		Or239280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239260_o0,
			i1 => And211940_o0,
			o0 => Or239280_o0
		);
		And239300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239280_o0,
			i1 => i12,
			o0 => And239300_o0
		);
		And239320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => Not180_o0,
			o0 => And239320_o0
		);
		And239340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => Nor22900_o0,
			o0 => And239340_o0
		);
		And239360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239340_o0,
			i1 => And239320_o0,
			o0 => And239360_o0
		);
		Or239380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239360_o0,
			i1 => And239300_o0,
			o0 => Or239380_o0
		);
		And239400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239380_o0,
			i1 => Not540_o0,
			o0 => And239400_o0
		);
		And239420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225680_o0,
			i1 => i12,
			o0 => And239420_o0
		);
		Or239440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239420_o0,
			i1 => And225060_o0,
			o0 => Or239440_o0
		);
		And239460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21060_o0,
			i1 => Not620_o0,
			o0 => And239460_o0
		);
		Or239480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239460_o0,
			i1 => And227220_o0,
			o0 => Or239480_o0
		);
		And239500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239480_o0,
			i1 => i5,
			o0 => And239500_o0
		);
		And239520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22900_o0,
			i1 => Nor21980_o0,
			o0 => And239520_o0
		);
		Or239540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239520_o0,
			i1 => And239500_o0,
			o0 => Or239540_o0
		);
		And239560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239540_o0,
			i1 => Or239440_o0,
			o0 => And239560_o0
		);
		And239580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => Not2080_o0,
			o0 => And239580_o0
		);
		And239600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239580_o0,
			i1 => Not180_o0,
			o0 => And239600_o0
		);
		And239620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1080_o0,
			i1 => i13,
			o0 => And239620_o0
		);
		And239640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239620_o0,
			i1 => i12,
			o0 => And239640_o0
		);
		Or239660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239640_o0,
			i1 => And239600_o0,
			o0 => Or239660_o0
		);
		And239680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239660_o0,
			i1 => And227220_o0,
			o0 => And239680_o0
		);
		And239700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239320_o0,
			i1 => And219800_o0,
			o0 => And239700_o0
		);
		Or239720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239700_o0,
			i1 => And239680_o0,
			o0 => Or239720_o0
		);
		And239740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239720_o0,
			i1 => i5,
			o0 => And239740_o0
		);
		And239760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => Not540_o0,
			o0 => And239760_o0
		);
		And239780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor224000_o0,
			i1 => i5,
			o0 => And239780_o0
		);
		Or239800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239780_o0,
			i1 => And239760_o0,
			o0 => Or239800_o0
		);
		And239820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239800_o0,
			i1 => And22800_o0,
			o0 => And239820_o0
		);
		And239840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239780_o0,
			i1 => And217280_o0,
			o0 => And239840_o0
		);
		And239860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225220_o0,
			i1 => And211020_o0,
			o0 => And239860_o0
		);
		And239880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239860_o0,
			i1 => And21120_o0,
			o0 => And239880_o0
		);
		Or239900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And239880_o0,
			i1 => And239840_o0,
			o0 => Or239900_o0
		);
		Or239920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239900_o0,
			i1 => And239820_o0,
			o0 => Or239920_o0
		);
		Or239940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239920_o0,
			i1 => And239740_o0,
			o0 => Or239940_o0
		);
		Or239960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239940_o0,
			i1 => And239560_o0,
			o0 => Or239960_o0
		);
		Or239980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239960_o0,
			i1 => And239400_o0,
			o0 => Or239980_o0
		);
		And240000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or239980_o0,
			i1 => And24040_o0,
			o0 => And240000_o0
		);
		Or240020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240000_o0,
			i1 => Nor233300_o0,
			o0 => Or240020_o0
		);
		And240040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230720_o0,
			i1 => Nor23600_o0,
			o0 => And240040_o0
		);
		And240060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240040_o0,
			i1 => Or240020_o0,
			o0 => And240060_o0
		);
		Or240080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240060_o0,
			i1 => And239200_o0,
			o0 => Or240080_o0
		);
		Or240100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or240080_o0,
			i1 => i36,
			o0 => Or240100_o0
		);
		And240120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240100_o0,
			i1 => And23700_o0,
			o0 => And240120_o0
		);
		And240140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i9,
			i1 => Not12100_o0,
			o0 => And240140_o0
		);
		And240160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => Not20520_o0,
			o0 => And240160_o0
		);
		And240180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240160_o0,
			i1 => Not12100_o0,
			o0 => And240180_o0
		);
		Or240200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240180_o0,
			i1 => And240140_o0,
			o0 => Or240200_o0
		);
		Or240220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or240200_o0,
			i1 => And235080_o0,
			o0 => Or240220_o0
		);
		Or240240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or240220_o0,
			i1 => And240120_o0,
			o0 => Or240240_o0
		);
		And240260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => i29,
			o0 => And240260_o0
		);
		And240280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240260_o0,
			i1 => And224320_o0,
			o0 => And240280_o0
		);
		Or240300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233720_o0,
			i1 => And218160_o0,
			o0 => Or240300_o0
		);
		And240320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i21,
			i1 => Not1500_o0,
			o0 => And240320_o0
		);
		And240340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240320_o0,
			i1 => And21640_o0,
			o0 => And240340_o0
		);
		And240360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i3,
			o0 => And240360_o0
		);
		And240380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240360_o0,
			i1 => Nor215260_o0,
			o0 => And240380_o0
		);
		And240400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240380_o0,
			i1 => And240340_o0,
			o0 => And240400_o0
		);
		And240420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240400_o0,
			i1 => Or240300_o0,
			o0 => And240420_o0
		);
		Or240440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240420_o0,
			i1 => And240280_o0,
			o0 => Or240440_o0
		);
		And240460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240440_o0,
			i1 => Not9540_o0,
			o0 => And240460_o0
		);
		And240480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i23,
			i1 => Not9800_o0,
			o0 => And240480_o0
		);
		Or240500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240480_o0,
			i1 => Not10520_o0,
			o0 => Or240500_o0
		);
		And240520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240500_o0,
			i1 => And240280_o0,
			o0 => And240520_o0
		);
		And240540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => Not1500_o0,
			o0 => And240540_o0
		);
		And240560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240380_o0,
			i1 => Nor218260_o0,
			o0 => And240560_o0
		);
		And240580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240560_o0,
			i1 => And240540_o0,
			o0 => And240580_o0
		);
		Or240600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240580_o0,
			i1 => And240520_o0,
			o0 => Or240600_o0
		);
		And240620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240600_o0,
			i1 => i20,
			o0 => And240620_o0
		);
		And240640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => Not32620_o0,
			o0 => And240640_o0
		);
		And240660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240640_o0,
			i1 => And224320_o0,
			o0 => And240660_o0
		);
		Or240680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240660_o0,
			i1 => And240620_o0,
			o0 => Or240680_o0
		);
		Or240700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or240680_o0,
			i1 => And240460_o0,
			o0 => Or240700_o0
		);
		And240720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240700_o0,
			i1 => i12,
			o0 => And240720_o0
		);
		And240740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i3,
			o0 => And240740_o0
		);
		Nor240760 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i3,
			o0 => Nor240760_o0
		);
		And240780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor240760_o0,
			i1 => And24940_o0,
			o0 => And240780_o0
		);
		Or240800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240780_o0,
			i1 => And240740_o0,
			o0 => Or240800_o0
		);
		And240820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240800_o0,
			i1 => i19,
			o0 => And240820_o0
		);
		And240840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor240760_o0,
			i1 => And222140_o0,
			o0 => And240840_o0
		);
		Or240860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240840_o0,
			i1 => And240820_o0,
			o0 => Or240860_o0
		);
		And240880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240860_o0,
			i1 => i17,
			o0 => And240880_o0
		);
		And240900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor236400_o0,
			i1 => Not140_o0,
			o0 => And240900_o0
		);
		And240920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240900_o0,
			i1 => And222140_o0,
			o0 => And240920_o0
		);
		Or240940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240920_o0,
			i1 => And240880_o0,
			o0 => Or240940_o0
		);
		And240960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240940_o0,
			i1 => And211340_o0,
			o0 => And240960_o0
		);
		Or240980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And240960_o0,
			i1 => And240720_o0,
			o0 => Or240980_o0
		);
		And241000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or240980_o0,
			i1 => Not620_o0,
			o0 => And241000_o0
		);
		Or241020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And222120_o0,
			i1 => i3,
			o0 => Or241020_o0
		);
		And241040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241020_o0,
			i1 => Nor2220_o0,
			o0 => And241040_o0
		);
		And241060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => i18,
			o0 => And241060_o0
		);
		And241080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241060_o0,
			i1 => And237940_o0,
			o0 => And241080_o0
		);
		Or241100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241080_o0,
			i1 => And241040_o0,
			o0 => Or241100_o0
		);
		And241120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241100_o0,
			i1 => Not1280_o0,
			o0 => And241120_o0
		);
		Or241140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => i3,
			o0 => Or241140_o0
		);
		And241160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21060_o0,
			i1 => Not1080_o0,
			o0 => And241160_o0
		);
		And241180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241160_o0,
			i1 => Or241140_o0,
			o0 => And241180_o0
		);
		Or241200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241180_o0,
			i1 => And241120_o0,
			o0 => Or241200_o0
		);
		And241220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241200_o0,
			i1 => Not540_o0,
			o0 => And241220_o0
		);
		And241240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor2960_o0,
			i1 => i3,
			o0 => And241240_o0
		);
		Or241260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241240_o0,
			i1 => Not7440_o0,
			o0 => Or241260_o0
		);
		And241280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i5,
			o0 => And241280_o0
		);
		And241300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241280_o0,
			i1 => Not1080_o0,
			o0 => And241300_o0
		);
		And241320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241300_o0,
			i1 => Or241260_o0,
			o0 => And241320_o0
		);
		Or241340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241320_o0,
			i1 => And241220_o0,
			o0 => Or241340_o0
		);
		And241360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => i15,
			o0 => And241360_o0
		);
		And241380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241360_o0,
			i1 => Or241340_o0,
			o0 => And241380_o0
		);
		Or241400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241380_o0,
			i1 => And241000_o0,
			o0 => Or241400_o0
		);
		And241420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241400_o0,
			i1 => Not120_o0,
			o0 => And241420_o0
		);
		And241440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			i1 => i18,
			o0 => And241440_o0
		);
		And241460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241440_o0,
			i1 => And22300_o0,
			o0 => And241460_o0
		);
		And241480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222820_o0,
			i1 => And23080_o0,
			o0 => And241480_o0
		);
		And241500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241480_o0,
			i1 => And241460_o0,
			o0 => And241500_o0
		);
		Or241520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241500_o0,
			i1 => And211160_o0,
			o0 => Or241520_o0
		);
		And241540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241520_o0,
			i1 => i5,
			o0 => And241540_o0
		);
		And241560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => Not620_o0,
			o0 => And241560_o0
		);
		And241580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29560_o0,
			i1 => And23080_o0,
			o0 => And241580_o0
		);
		And241600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241580_o0,
			i1 => And233960_o0,
			o0 => And241600_o0
		);
		And241620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241600_o0,
			i1 => And241560_o0,
			o0 => And241620_o0
		);
		Or241640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241620_o0,
			i1 => And211160_o0,
			o0 => Or241640_o0
		);
		And241660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241640_o0,
			i1 => Not540_o0,
			o0 => And241660_o0
		);
		Or241680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241660_o0,
			i1 => And241540_o0,
			o0 => Or241680_o0
		);
		And241700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241680_o0,
			i1 => Not1500_o0,
			o0 => And241700_o0
		);
		And241720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And241360_o0,
			i1 => And218580_o0,
			o0 => And241720_o0
		);
		Or241740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241720_o0,
			i1 => And241700_o0,
			o0 => Or241740_o0
		);
		And241760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241740_o0,
			i1 => Not1280_o0,
			o0 => And241760_o0
		);
		Or241780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241760_o0,
			i1 => And211360_o0,
			o0 => Or241780_o0
		);
		And241800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241780_o0,
			i1 => Not140_o0,
			o0 => And241800_o0
		);
		Or241820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241800_o0,
			i1 => And211480_o0,
			o0 => Or241820_o0
		);
		And241840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241820_o0,
			i1 => i2,
			o0 => And241840_o0
		);
		Or241860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241840_o0,
			i1 => And241420_o0,
			o0 => Or241860_o0
		);
		And241880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241860_o0,
			i1 => Not160_o0,
			o0 => And241880_o0
		);
		And241900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211460_o0,
			i1 => i4,
			o0 => And241900_o0
		);
		Or241920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241900_o0,
			i1 => And241880_o0,
			o0 => Or241920_o0
		);
		And241940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241920_o0,
			i1 => Not100_o0,
			o0 => And241940_o0
		);
		Or241960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And241940_o0,
			i1 => And211620_o0,
			o0 => Or241960_o0
		);
		And241980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or241960_o0,
			i1 => Not60_o0,
			o0 => And241980_o0
		);
		And242000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or231100_o0,
			i1 => And23020_o0,
			o0 => And242000_o0
		);
		And242020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23180_o0,
			i1 => Not120_o0,
			o0 => And242020_o0
		);
		And242040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242020_o0,
			i1 => And242000_o0,
			o0 => And242040_o0
		);
		Or242060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242040_o0,
			i1 => And241980_o0,
			o0 => Or242060_o0
		);
		And242080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242060_o0,
			i1 => Not80_o0,
			o0 => And242080_o0
		);
		And242100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => Nor21140_o0,
			o0 => And242100_o0
		);
		And242120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242100_o0,
			i1 => Nor23600_o0,
			o0 => And242120_o0
		);
		Or242140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i15,
			o0 => Or242140_o0
		);
		And242160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And226340_o0,
			i1 => And212000_o0,
			o0 => And242160_o0
		);
		And242180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242160_o0,
			i1 => Or242140_o0,
			o0 => And242180_o0
		);
		And242200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242180_o0,
			i1 => And242120_o0,
			o0 => And242200_o0
		);
		Or242220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242200_o0,
			i1 => And242080_o0,
			o0 => Or242220_o0
		);
		And242240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242220_o0,
			i1 => And23360_o0,
			o0 => And242240_o0
		);
		And242260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i2,
			o0 => And242260_o0
		);
		And242280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242260_o0,
			i1 => And230320_o0,
			o0 => And242280_o0
		);
		And242300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24940_o0,
			i1 => Not120_o0,
			o0 => And242300_o0
		);
		Or242320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242300_o0,
			i1 => And242280_o0,
			o0 => Or242320_o0
		);
		And242340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242320_o0,
			i1 => Nor240760_o0,
			o0 => And242340_o0
		);
		And242360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i5,
			o0 => And242360_o0
		);
		And242380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242360_o0,
			i1 => And26040_o0,
			o0 => And242380_o0
		);
		And242400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242380_o0,
			i1 => Or229560_o0,
			o0 => And242400_o0
		);
		Or242420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242400_o0,
			i1 => And242340_o0,
			o0 => Or242420_o0
		);
		And242440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242420_o0,
			i1 => And22300_o0,
			o0 => And242440_o0
		);
		And242460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor240760_o0,
			i1 => Not120_o0,
			o0 => And242460_o0
		);
		And242480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24180_o0,
			i1 => And22800_o0,
			o0 => And242480_o0
		);
		And242500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242480_o0,
			i1 => And242460_o0,
			o0 => And242500_o0
		);
		Or242520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242500_o0,
			i1 => And242440_o0,
			o0 => Or242520_o0
		);
		And242540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242520_o0,
			i1 => And23080_o0,
			o0 => And242540_o0
		);
		And242560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210400_o0,
			i1 => Not140_o0,
			o0 => And242560_o0
		);
		And242580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242560_o0,
			i1 => Not120_o0,
			o0 => And242580_o0
		);
		Or242600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242580_o0,
			i1 => Or23980_o0,
			o0 => Or242600_o0
		);
		And242620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And27500_o0,
			i1 => And23020_o0,
			o0 => And242620_o0
		);
		And242640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242620_o0,
			i1 => Or242600_o0,
			o0 => And242640_o0
		);
		Or242660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242640_o0,
			i1 => And242540_o0,
			o0 => Or242660_o0
		);
		And242680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242660_o0,
			i1 => Not1280_o0,
			o0 => And242680_o0
		);
		Or242700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or210400_o0,
			i1 => i3,
			o0 => Or242700_o0
		);
		And242720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242700_o0,
			i1 => i15,
			o0 => And242720_o0
		);
		And242740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor240760_o0,
			i1 => And223380_o0,
			o0 => And242740_o0
		);
		Or242760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242740_o0,
			i1 => And242720_o0,
			o0 => Or242760_o0
		);
		And242780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242760_o0,
			i1 => Not1040_o0,
			o0 => And242780_o0
		);
		And242800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223240_o0,
			i1 => Not620_o0,
			o0 => And242800_o0
		);
		And242820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242800_o0,
			i1 => Nor240760_o0,
			o0 => And242820_o0
		);
		Or242840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242820_o0,
			i1 => And242780_o0,
			o0 => Or242840_o0
		);
		And242860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242840_o0,
			i1 => And23020_o0,
			o0 => And242860_o0
		);
		And242880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210020_o0,
			i1 => And22300_o0,
			o0 => And242880_o0
		);
		Or242900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242880_o0,
			i1 => i15,
			o0 => Or242900_o0
		);
		And242920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => i40,
			o0 => And242920_o0
		);
		And242940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242920_o0,
			i1 => Nor240760_o0,
			o0 => And242940_o0
		);
		And242960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And242940_o0,
			i1 => Or242900_o0,
			o0 => And242960_o0
		);
		Or242980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242960_o0,
			i1 => And242860_o0,
			o0 => Or242980_o0
		);
		And243000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or242980_o0,
			i1 => Not1080_o0,
			o0 => And243000_o0
		);
		And243020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24180_o0,
			i1 => And23080_o0,
			o0 => And243020_o0
		);
		And243040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243020_o0,
			i1 => Nor240760_o0,
			o0 => And243040_o0
		);
		And243060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243040_o0,
			i1 => Or231500_o0,
			o0 => And243060_o0
		);
		Or243080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243060_o0,
			i1 => And243000_o0,
			o0 => Or243080_o0
		);
		And243100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243080_o0,
			i1 => Not120_o0,
			o0 => And243100_o0
		);
		And243120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211160_o0,
			i1 => i2,
			o0 => And243120_o0
		);
		Or243140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243120_o0,
			i1 => And243100_o0,
			o0 => Or243140_o0
		);
		And243160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243140_o0,
			i1 => i16,
			o0 => And243160_o0
		);
		Or243180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243160_o0,
			i1 => And242680_o0,
			o0 => Or243180_o0
		);
		And243200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243180_o0,
			i1 => Not1500_o0,
			o0 => And243200_o0
		);
		And243220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223960_o0,
			i1 => And215820_o0,
			o0 => And243220_o0
		);
		Or243240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243220_o0,
			i1 => Not1280_o0,
			o0 => Or243240_o0
		);
		And243260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243240_o0,
			i1 => Not180_o0,
			o0 => And243260_o0
		);
		Or243280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i23,
			i1 => i22,
			o0 => Or243280_o0
		);
		And243300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			i1 => i12,
			o0 => And243300_o0
		);
		And243320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i29,
			i1 => i21,
			o0 => And243320_o0
		);
		And243340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243320_o0,
			i1 => And243300_o0,
			o0 => And243340_o0
		);
		And243360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243340_o0,
			i1 => Or243280_o0,
			o0 => And243360_o0
		);
		Or243380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243360_o0,
			i1 => And243260_o0,
			o0 => Or243380_o0
		);
		And243400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243380_o0,
			i1 => Not620_o0,
			o0 => And243400_o0
		);
		Nor243420 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor26980_o0,
			i1 => i16,
			o0 => Nor243420_o0
		);
		Or243440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor243420_o0,
			i1 => And2320_o0,
			o0 => Or243440_o0
		);
		And243460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233000_o0,
			i1 => i19,
			o0 => And243460_o0
		);
		And243480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243460_o0,
			i1 => Or243440_o0,
			o0 => And243480_o0
		);
		Or243500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243480_o0,
			i1 => And243400_o0,
			o0 => Or243500_o0
		);
		And243520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243500_o0,
			i1 => And2560_o0,
			o0 => And243520_o0
		);
		And243540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210940_o0,
			i1 => Not180_o0,
			o0 => And243540_o0
		);
		And243560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243540_o0,
			i1 => i5,
			o0 => And243560_o0
		);
		Or243580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243560_o0,
			i1 => And243520_o0,
			o0 => Or243580_o0
		);
		And243600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243580_o0,
			i1 => Not140_o0,
			o0 => And243600_o0
		);
		And243620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243540_o0,
			i1 => i3,
			o0 => And243620_o0
		);
		Or243640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243620_o0,
			i1 => And243600_o0,
			o0 => Or243640_o0
		);
		And243660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243640_o0,
			i1 => Not120_o0,
			o0 => And243660_o0
		);
		And243680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243540_o0,
			i1 => i2,
			o0 => And243680_o0
		);
		Or243700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243680_o0,
			i1 => And243660_o0,
			o0 => Or243700_o0
		);
		And243720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243700_o0,
			i1 => i13,
			o0 => And243720_o0
		);
		Or243740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not1040_o0,
			i1 => i16,
			o0 => Or243740_o0
		);
		Or243760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or243740_o0,
			i1 => And219940_o0,
			o0 => Or243760_o0
		);
		And243780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243760_o0,
			i1 => i15,
			o0 => And243780_o0
		);
		Or243800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243780_o0,
			i1 => And227280_o0,
			o0 => Or243800_o0
		);
		And243820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not2080_o0,
			o0 => And243820_o0
		);
		And243840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243820_o0,
			i1 => Nor21140_o0,
			o0 => And243840_o0
		);
		And243860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243840_o0,
			i1 => And236920_o0,
			o0 => And243860_o0
		);
		And243880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243860_o0,
			i1 => Or243800_o0,
			o0 => And243880_o0
		);
		Or243900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And243880_o0,
			i1 => And243720_o0,
			o0 => Or243900_o0
		);
		Or243920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or243900_o0,
			i1 => And243200_o0,
			o0 => Or243920_o0
		);
		And243940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or243920_o0,
			i1 => Not160_o0,
			o0 => And243940_o0
		);
		And243960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240360_o0,
			i1 => Not120_o0,
			o0 => And243960_o0
		);
		And243980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243960_o0,
			i1 => And230540_o0,
			o0 => And243980_o0
		);
		And244000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And243980_o0,
			i1 => And230520_o0,
			o0 => And244000_o0
		);
		Or244020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244000_o0,
			i1 => And211460_o0,
			o0 => Or244020_o0
		);
		And244040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244020_o0,
			i1 => i4,
			o0 => And244040_o0
		);
		Or244060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244040_o0,
			i1 => And243940_o0,
			o0 => Or244060_o0
		);
		And244080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244060_o0,
			i1 => Not100_o0,
			o0 => And244080_o0
		);
		Or244100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244080_o0,
			i1 => And211620_o0,
			o0 => Or244100_o0
		);
		And244120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244100_o0,
			i1 => Not80_o0,
			o0 => And244120_o0
		);
		And244140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225460_o0,
			i1 => Nor215260_o0,
			o0 => And244140_o0
		);
		Or244160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244140_o0,
			i1 => i13,
			o0 => Or244160_o0
		);
		And244180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244160_o0,
			i1 => Not180_o0,
			o0 => And244180_o0
		);
		Or244200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => And216160_o0,
			o0 => Or244200_o0
		);
		And244220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244200_o0,
			i1 => Not1280_o0,
			o0 => And244220_o0
		);
		Or244240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244220_o0,
			i1 => And21120_o0,
			o0 => Or244240_o0
		);
		Or244260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244240_o0,
			i1 => Not2080_o0,
			o0 => Or244260_o0
		);
		And244280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244260_o0,
			i1 => i12,
			o0 => And244280_o0
		);
		Or244300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244280_o0,
			i1 => And244180_o0,
			o0 => Or244300_o0
		);
		And244320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244300_o0,
			i1 => Not620_o0,
			o0 => And244320_o0
		);
		And244340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => i17,
			o0 => And244340_o0
		);
		And244360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor238120_o0,
			i1 => Not180_o0,
			o0 => And244360_o0
		);
		Or244380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244360_o0,
			i1 => And244340_o0,
			o0 => Or244380_o0
		);
		And244400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244380_o0,
			i1 => And2640_o0,
			o0 => And244400_o0
		);
		And244420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225240_o0,
			i1 => And219800_o0,
			o0 => And244420_o0
		);
		Or244440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i15,
			o0 => Or244440_o0
		);
		And244460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244440_o0,
			i1 => Nor224000_o0,
			o0 => And244460_o0
		);
		And244480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228580_o0,
			i1 => And28120_o0,
			o0 => And244480_o0
		);
		Or244500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244480_o0,
			i1 => And244460_o0,
			o0 => Or244500_o0
		);
		Or244520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244500_o0,
			i1 => And244420_o0,
			o0 => Or244520_o0
		);
		Or244540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244520_o0,
			i1 => And244400_o0,
			o0 => Or244540_o0
		);
		Or244560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244540_o0,
			i1 => And244320_o0,
			o0 => Or244560_o0
		);
		And244580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217680_o0,
			i1 => And22620_o0,
			o0 => And244580_o0
		);
		And244600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And244580_o0,
			i1 => Or244560_o0,
			o0 => And244600_o0
		);
		Or244620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244600_o0,
			i1 => And244120_o0,
			o0 => Or244620_o0
		);
		And244640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244620_o0,
			i1 => Not60_o0,
			o0 => And244640_o0
		);
		And244660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => And28900_o0,
			o0 => And244660_o0
		);
		Or244680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244660_o0,
			i1 => And28860_o0,
			o0 => Or244680_o0
		);
		And244700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244680_o0,
			i1 => i16,
			o0 => And244700_o0
		);
		Or244720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244700_o0,
			i1 => And231060_o0,
			o0 => Or244720_o0
		);
		And244740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244720_o0,
			i1 => And224880_o0,
			o0 => And244740_o0
		);
		Or244760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244740_o0,
			i1 => And244640_o0,
			o0 => Or244760_o0
		);
		And244780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244760_o0,
			i1 => And23360_o0,
			o0 => And244780_o0
		);
		And244800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i24,
			o0 => And244800_o0
		);
		And244820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			i1 => Not9540_o0,
			o0 => And244820_o0
		);
		And244840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And244820_o0,
			i1 => i23,
			o0 => And244840_o0
		);
		And244860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And244840_o0,
			i1 => And244800_o0,
			o0 => And244860_o0
		);
		Or244880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244860_o0,
			i1 => i20,
			o0 => Or244880_o0
		);
		And244900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244880_o0,
			i1 => And240320_o0,
			o0 => And244900_o0
		);
		Or244920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244900_o0,
			i1 => i19,
			o0 => Or244920_o0
		);
		Or244940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244920_o0,
			i1 => Not1080_o0,
			o0 => Or244940_o0
		);
		Or244960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244940_o0,
			i1 => i16,
			o0 => Or244960_o0
		);
		Or244980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or244960_o0,
			i1 => Not1040_o0,
			o0 => Or244980_o0
		);
		And245000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244980_o0,
			i1 => Not2080_o0,
			o0 => And245000_o0
		);
		Or245020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217800_o0,
			i1 => Nand210560_o0,
			o0 => Or245020_o0
		);
		And245040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245020_o0,
			i1 => And29560_o0,
			o0 => And245040_o0
		);
		Or245060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245040_o0,
			i1 => And210540_o0,
			o0 => Or245060_o0
		);
		And245080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240540_o0,
			i1 => Nor215260_o0,
			o0 => And245080_o0
		);
		And245100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245080_o0,
			i1 => Or245060_o0,
			o0 => And245100_o0
		);
		And245120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => i13,
			o0 => And245120_o0
		);
		And245140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245120_o0,
			i1 => And2400_o0,
			o0 => And245140_o0
		);
		Or245160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245140_o0,
			i1 => And245100_o0,
			o0 => Or245160_o0
		);
		And245180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29720_o0,
			i1 => i23,
			o0 => And245180_o0
		);
		And245200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245180_o0,
			i1 => Nor215260_o0,
			o0 => And245200_o0
		);
		And245220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234540_o0,
			i1 => Not9540_o0,
			o0 => And245220_o0
		);
		And245240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245220_o0,
			i1 => And228740_o0,
			o0 => And245240_o0
		);
		And245260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245240_o0,
			i1 => And245200_o0,
			o0 => And245260_o0
		);
		And245280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not7120_o0,
			i1 => i13,
			o0 => And245280_o0
		);
		And245300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245280_o0,
			i1 => i28,
			o0 => And245300_o0
		);
		Or245320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245300_o0,
			i1 => And245260_o0,
			o0 => Or245320_o0
		);
		And245340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not7140_o0,
			i1 => i24,
			o0 => And245340_o0
		);
		Or245360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245340_o0,
			i1 => Not3840_o0,
			o0 => Or245360_o0
		);
		And245380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245360_o0,
			i1 => i13,
			o0 => And245380_o0
		);
		Or245400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245380_o0,
			i1 => Or245320_o0,
			o0 => Or245400_o0
		);
		Or245420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or245400_o0,
			i1 => Or245160_o0,
			o0 => Or245420_o0
		);
		Or245440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or245420_o0,
			i1 => And245000_o0,
			o0 => Or245440_o0
		);
		And245460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245440_o0,
			i1 => i12,
			o0 => And245460_o0
		);
		Or245480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or219240_o0,
			i1 => And23440_o0,
			o0 => Or245480_o0
		);
		And245500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245480_o0,
			i1 => Not180_o0,
			o0 => And245500_o0
		);
		Or245520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245500_o0,
			i1 => And245460_o0,
			o0 => Or245520_o0
		);
		And245540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245520_o0,
			i1 => Not620_o0,
			o0 => And245540_o0
		);
		Nand245560 : entity gtech_lib.nand2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => Not12240_o0,
			o0 => Nand245560_o0
		);
		Or245580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand245560_o0,
			i1 => i19,
			o0 => Or245580_o0
		);
		And245600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215260_o0,
			i1 => Nor2220_o0,
			o0 => And245600_o0
		);
		And245620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And245600_o0,
			i1 => Or245580_o0,
			o0 => And245620_o0
		);
		Or245640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245620_o0,
			i1 => i13,
			o0 => Or245640_o0
		);
		And245660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245640_o0,
			i1 => i12,
			o0 => And245660_o0
		);
		Xor245680 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => i12,
			o0 => Xor245680_o0
		);
		And245700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor245680_o0,
			i1 => And21940_o0,
			o0 => And245700_o0
		);
		And245720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219240_o0,
			i1 => Not180_o0,
			o0 => And245720_o0
		);
		And245740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => i16,
			o0 => And245740_o0
		);
		Or245760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245740_o0,
			i1 => And245720_o0,
			o0 => Or245760_o0
		);
		Or245780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or245760_o0,
			i1 => And245700_o0,
			o0 => Or245780_o0
		);
		Or245800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand245560_o0,
			i1 => Not1080_o0,
			o0 => Or245800_o0
		);
		And245820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245800_o0,
			i1 => And23020_o0,
			o0 => And245820_o0
		);
		And245840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239580_o0,
			i1 => i12,
			o0 => And245840_o0
		);
		Or245860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245840_o0,
			i1 => And245820_o0,
			o0 => Or245860_o0
		);
		And245880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245860_o0,
			i1 => Nor22900_o0,
			o0 => And245880_o0
		);
		Or245900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245880_o0,
			i1 => Or245780_o0,
			o0 => Or245900_o0
		);
		Or245920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or245900_o0,
			i1 => And245660_o0,
			o0 => Or245920_o0
		);
		And245940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245920_o0,
			i1 => i15,
			o0 => And245940_o0
		);
		Or245960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And245940_o0,
			i1 => And245540_o0,
			o0 => Or245960_o0
		);
		And245980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or245960_o0,
			i1 => Not80_o0,
			o0 => And245980_o0
		);
		Xor246000 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => i12,
			o0 => Xor246000_o0
		);
		Not46020 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Xor246000_o0,
			o0 => Not46020_o0
		);
		Or246040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not46020_o0,
			i1 => Xor245680_o0,
			o0 => Or246040_o0
		);
		And246060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246040_o0,
			i1 => i14,
			o0 => And246060_o0
		);
		Or246080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246060_o0,
			i1 => And245980_o0,
			o0 => Or246080_o0
		);
		Or246100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or246080_o0,
			i1 => Not24560_o0,
			o0 => Or246100_o0
		);
		And246120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246100_o0,
			i1 => Nor214960_o0,
			o0 => And246120_o0
		);
		Or246140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246120_o0,
			i1 => i8,
			o0 => Or246140_o0
		);
		And246160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246140_o0,
			i1 => Not540_o0,
			o0 => And246160_o0
		);
		And246180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24040_o0,
			i1 => Not180_o0,
			o0 => And246180_o0
		);
		And246200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231400_o0,
			i1 => And213900_o0,
			o0 => And246200_o0
		);
		Or246220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246200_o0,
			i1 => And246180_o0,
			o0 => Or246220_o0
		);
		And246240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246220_o0,
			i1 => Not620_o0,
			o0 => And246240_o0
		);
		And246260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not80_o0,
			o0 => And246260_o0
		);
		And246280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246260_o0,
			i1 => i12,
			o0 => And246280_o0
		);
		Or246300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246280_o0,
			i1 => And227100_o0,
			o0 => Or246300_o0
		);
		And246320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i15,
			o0 => And246320_o0
		);
		And246340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246320_o0,
			i1 => Or246300_o0,
			o0 => And246340_o0
		);
		Or246360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246340_o0,
			i1 => And246240_o0,
			o0 => Or246360_o0
		);
		And246380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246360_o0,
			i1 => Not1280_o0,
			o0 => And246380_o0
		);
		And246400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => i12,
			o0 => And246400_o0
		);
		Or246420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246400_o0,
			i1 => And227100_o0,
			o0 => Or246420_o0
		);
		And246440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246420_o0,
			i1 => And28480_o0,
			o0 => And246440_o0
		);
		Or246460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246440_o0,
			i1 => And246380_o0,
			o0 => Or246460_o0
		);
		And246480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246460_o0,
			i1 => i18,
			o0 => And246480_o0
		);
		Or246500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227100_o0,
			i1 => And227060_o0,
			o0 => Or246500_o0
		);
		And246520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246500_o0,
			i1 => i40,
			o0 => And246520_o0
		);
		And246540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228340_o0,
			i1 => And213900_o0,
			o0 => And246540_o0
		);
		Or246560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246540_o0,
			i1 => And246520_o0,
			o0 => Or246560_o0
		);
		And246580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246560_o0,
			i1 => Not1080_o0,
			o0 => And246580_o0
		);
		Or246600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246580_o0,
			i1 => And246480_o0,
			o0 => Or246600_o0
		);
		And246620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246600_o0,
			i1 => i17,
			o0 => And246620_o0
		);
		And246640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or227080_o0,
			i1 => i40,
			o0 => And246640_o0
		);
		And246660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2240_o0,
			i1 => Not1280_o0,
			o0 => And246660_o0
		);
		And246680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246660_o0,
			i1 => And246400_o0,
			o0 => And246680_o0
		);
		Or246700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246680_o0,
			i1 => And246640_o0,
			o0 => Or246700_o0
		);
		And246720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246700_o0,
			i1 => Not1040_o0,
			o0 => And246720_o0
		);
		Or246740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246720_o0,
			i1 => And246620_o0,
			o0 => Or246740_o0
		);
		And246760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or246740_o0,
			i1 => Not2080_o0,
			o0 => And246760_o0
		);
		And246780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not28160_o0,
			i1 => And2640_o0,
			o0 => And246780_o0
		);
		And246800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => And21300_o0,
			o0 => And246800_o0
		);
		Or246820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246800_o0,
			i1 => And246780_o0,
			o0 => Or246820_o0
		);
		And246840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24000_o0,
			i1 => i17,
			o0 => And246840_o0
		);
		And246860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246840_o0,
			i1 => Or246820_o0,
			o0 => And246860_o0
		);
		Or246880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And24620_o0,
			i1 => i15,
			o0 => Or246880_o0
		);
		And246900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223240_o0,
			i1 => And22560_o0,
			o0 => And246900_o0
		);
		And246920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246900_o0,
			i1 => Or246880_o0,
			o0 => And246920_o0
		);
		And246940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212220_o0,
			i1 => Nor24000_o0,
			o0 => And246940_o0
		);
		And246960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => i12,
			o0 => And246960_o0
		);
		And246980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246960_o0,
			i1 => And216040_o0,
			o0 => And246980_o0
		);
		Or247000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And246980_o0,
			i1 => And246940_o0,
			o0 => Or247000_o0
		);
		And247020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => Not180_o0,
			o0 => And247020_o0
		);
		And247040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247020_o0,
			i1 => And2320_o0,
			o0 => And247040_o0
		);
		And247060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => And22560_o0,
			o0 => And247060_o0
		);
		And247080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247060_o0,
			i1 => And28280_o0,
			o0 => And247080_o0
		);
		Or247100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247080_o0,
			i1 => And247040_o0,
			o0 => Or247100_o0
		);
		Or247120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or247100_o0,
			i1 => Or247000_o0,
			o0 => Or247120_o0
		);
		Or247140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or247120_o0,
			i1 => And246920_o0,
			o0 => Or247140_o0
		);
		Or247160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or247140_o0,
			i1 => And246860_o0,
			o0 => Or247160_o0
		);
		And247180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247160_o0,
			i1 => i13,
			o0 => And247180_o0
		);
		Or247200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247180_o0,
			i1 => And246760_o0,
			o0 => Or247200_o0
		);
		And247220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227400_o0,
			i1 => Not12120_o0,
			o0 => And247220_o0
		);
		And247240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247220_o0,
			i1 => Or247200_o0,
			o0 => And247240_o0
		);
		Or247260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247240_o0,
			i1 => And246160_o0,
			o0 => Or247260_o0
		);
		And247280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247260_o0,
			i1 => Not160_o0,
			o0 => And247280_o0
		);
		And247300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or221040_o0,
			i1 => And211240_o0,
			o0 => And247300_o0
		);
		Or247320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247300_o0,
			i1 => And233660_o0,
			o0 => Or247320_o0
		);
		And247340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247320_o0,
			i1 => Not1500_o0,
			o0 => And247340_o0
		);
		Or247360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247340_o0,
			i1 => And237220_o0,
			o0 => Or247360_o0
		);
		And247380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247360_o0,
			i1 => i17,
			o0 => And247380_o0
		);
		And247400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239620_o0,
			i1 => Not180_o0,
			o0 => And247400_o0
		);
		And247420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => And2240_o0,
			o0 => And247420_o0
		);
		Or247440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247420_o0,
			i1 => And247400_o0,
			o0 => Or247440_o0
		);
		And247460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247440_o0,
			i1 => And22800_o0,
			o0 => And247460_o0
		);
		Or247480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247460_o0,
			i1 => And247380_o0,
			o0 => Or247480_o0
		);
		And247500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247480_o0,
			i1 => Not1280_o0,
			o0 => And247500_o0
		);
		Or247520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247500_o0,
			i1 => And211360_o0,
			o0 => Or247520_o0
		);
		And247540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247520_o0,
			i1 => Not80_o0,
			o0 => And247540_o0
		);
		And247560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12100_o0,
			i1 => i4,
			o0 => And247560_o0
		);
		And247580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247560_o0,
			i1 => Not12120_o0,
			o0 => And247580_o0
		);
		And247600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247580_o0,
			i1 => And247540_o0,
			o0 => And247600_o0
		);
		Or247620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247600_o0,
			i1 => And247280_o0,
			o0 => Or247620_o0
		);
		And247640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247620_o0,
			i1 => Not140_o0,
			o0 => And247640_o0
		);
		And247660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And238360_o0,
			i1 => Or217980_o0,
			o0 => And247660_o0
		);
		Nor247680 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => i4,
			o0 => Nor247680_o0
		);
		Or247700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor247680_o0,
			i1 => And247660_o0,
			o0 => Or247700_o0
		);
		And247720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247700_o0,
			i1 => And211240_o0,
			o0 => And247720_o0
		);
		And247740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233660_o0,
			i1 => Not160_o0,
			o0 => And247740_o0
		);
		Or247760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247740_o0,
			i1 => And247720_o0,
			o0 => Or247760_o0
		);
		And247780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247760_o0,
			i1 => Not1500_o0,
			o0 => And247780_o0
		);
		And247800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => Not160_o0,
			o0 => And247800_o0
		);
		And247820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247800_o0,
			i1 => And237200_o0,
			o0 => And247820_o0
		);
		Or247840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247820_o0,
			i1 => And247780_o0,
			o0 => Or247840_o0
		);
		And247860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247840_o0,
			i1 => And237260_o0,
			o0 => And247860_o0
		);
		Not47880 : entity gtech_lib.not_d
		generic map(1000 fs)
		port map(
			i0 => Nand210560_o0,
			o0 => Not47880_o0
		);
		Nor247900 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor218020_o0,
			i1 => Not47880_o0,
			o0 => Nor247900_o0
		);
		Or247920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor247900_o0,
			i1 => And221280_o0,
			o0 => Or247920_o0
		);
		And247940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247920_o0,
			i1 => And29560_o0,
			o0 => And247940_o0
		);
		Or247960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And247940_o0,
			i1 => And218280_o0,
			o0 => Or247960_o0
		);
		And247980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or247960_o0,
			i1 => Not1500_o0,
			o0 => And247980_o0
		);
		And248000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => And21640_o0,
			o0 => And248000_o0
		);
		And248020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248000_o0,
			i1 => And22100_o0,
			o0 => And248020_o0
		);
		And248040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248020_o0,
			i1 => And247980_o0,
			o0 => And248040_o0
		);
		Or248060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248040_o0,
			i1 => Or211280_o0,
			o0 => Or248060_o0
		);
		And248080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248060_o0,
			i1 => Not1280_o0,
			o0 => And248080_o0
		);
		Or248100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248080_o0,
			i1 => And211360_o0,
			o0 => Or248100_o0
		);
		Or248120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or248100_o0,
			i1 => And247860_o0,
			o0 => Or248120_o0
		);
		And248140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248120_o0,
			i1 => Not80_o0,
			o0 => And248140_o0
		);
		And248160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12100_o0,
			i1 => i3,
			o0 => And248160_o0
		);
		And248180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248160_o0,
			i1 => Not12120_o0,
			o0 => And248180_o0
		);
		And248200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248180_o0,
			i1 => And248140_o0,
			o0 => And248200_o0
		);
		Or248220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248200_o0,
			i1 => And247640_o0,
			o0 => Or248220_o0
		);
		And248240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248220_o0,
			i1 => Not120_o0,
			o0 => And248240_o0
		);
		And248260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => And29560_o0,
			o0 => And248260_o0
		);
		And248280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => And21940_o0,
			o0 => And248280_o0
		);
		And248300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222800_o0,
			i1 => Nor22600_o0,
			o0 => And248300_o0
		);
		And248320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248300_o0,
			i1 => And248280_o0,
			o0 => And248320_o0
		);
		And248340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248320_o0,
			i1 => And248260_o0,
			o0 => And248340_o0
		);
		And248360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248340_o0,
			i1 => And221460_o0,
			o0 => And248360_o0
		);
		Or248380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248360_o0,
			i1 => Or230440_o0,
			o0 => Or248380_o0
		);
		And248400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248380_o0,
			i1 => Not80_o0,
			o0 => And248400_o0
		);
		And248420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12100_o0,
			i1 => i2,
			o0 => And248420_o0
		);
		And248440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248420_o0,
			i1 => Not12120_o0,
			o0 => And248440_o0
		);
		And248460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248440_o0,
			i1 => And248400_o0,
			o0 => And248460_o0
		);
		Or248480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248460_o0,
			i1 => And248240_o0,
			o0 => Or248480_o0
		);
		And248500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248480_o0,
			i1 => Not100_o0,
			o0 => And248500_o0
		);
		And248520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not12100_o0,
			i1 => i1,
			o0 => And248520_o0
		);
		And248540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248520_o0,
			i1 => Not12120_o0,
			o0 => And248540_o0
		);
		And248560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248540_o0,
			i1 => And230860_o0,
			o0 => And248560_o0
		);
		Or248580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248560_o0,
			i1 => And248500_o0,
			o0 => Or248580_o0
		);
		And248600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248580_o0,
			i1 => Not60_o0,
			o0 => And248600_o0
		);
		Or248620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And242000_o0,
			i1 => And23140_o0,
			o0 => Or248620_o0
		);
		And248640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248620_o0,
			i1 => Not80_o0,
			o0 => And248640_o0
		);
		Nor248660 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i8,
			i1 => i2,
			o0 => Nor248660_o0
		);
		And248680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor248660_o0,
			i1 => Not12120_o0,
			o0 => And248680_o0
		);
		And248700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248680_o0,
			i1 => And23180_o0,
			o0 => And248700_o0
		);
		And248720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248700_o0,
			i1 => And248640_o0,
			o0 => And248720_o0
		);
		Or248740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248720_o0,
			i1 => And248600_o0,
			o0 => Or248740_o0
		);
		And248760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248740_o0,
			i1 => Not3300_o0,
			o0 => And248760_o0
		);
		Or248780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i10,
			o0 => Or248780_o0
		);
		And248800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248780_o0,
			i1 => Not12100_o0,
			o0 => And248800_o0
		);
		Or248820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248800_o0,
			i1 => And248760_o0,
			o0 => Or248820_o0
		);
		And248840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248820_o0,
			i1 => Not24960_o0,
			o0 => And248840_o0
		);
		And248860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or220620_o0,
			i1 => i11,
			o0 => And248860_o0
		);
		Or248880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248860_o0,
			i1 => And248840_o0,
			o0 => Or248880_o0
		);
		And248900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or248880_o0,
			i1 => Not20520_o0,
			o0 => And248900_o0
		);
		And248920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not24960_o0,
			i1 => i10,
			o0 => And248920_o0
		);
		And248940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248920_o0,
			i1 => And240140_o0,
			o0 => And248940_o0
		);
		Or248960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And248940_o0,
			i1 => And248900_o0,
			o0 => Or248960_o0
		);
		And248980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220200_o0,
			i1 => And213240_o0,
			o0 => And248980_o0
		);
		And249000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248980_o0,
			i1 => And212280_o0,
			o0 => And249000_o0
		);
		And249020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And249000_o0,
			i1 => Or225740_o0,
			o0 => And249020_o0
		);
		And249040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And249020_o0,
			i1 => And23640_o0,
			o0 => And249040_o0
		);
		Or249060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249040_o0,
			i1 => i10,
			o0 => Or249060_o0
		);
		And249080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249060_o0,
			i1 => Not20520_o0,
			o0 => And249080_o0
		);
		Or249100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249080_o0,
			i1 => And212160_o0,
			o0 => Or249100_o0
		);
		And249120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249100_o0,
			i1 => Not12100_o0,
			o0 => And249120_o0
		);
		Or249140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or220920_o0,
			i1 => Not1080_o0,
			o0 => Or249140_o0
		);
		And249160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249140_o0,
			i1 => And211240_o0,
			o0 => And249160_o0
		);
		Or249180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249160_o0,
			i1 => And233660_o0,
			o0 => Or249180_o0
		);
		And249200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249180_o0,
			i1 => Not1500_o0,
			o0 => And249200_o0
		);
		Or249220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249200_o0,
			i1 => And237220_o0,
			o0 => Or249220_o0
		);
		And249240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249220_o0,
			i1 => i17,
			o0 => And249240_o0
		);
		Or249260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249240_o0,
			i1 => And247460_o0,
			o0 => Or249260_o0
		);
		And249280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249260_o0,
			i1 => Not1280_o0,
			o0 => And249280_o0
		);
		And249300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229800_o0,
			i1 => And23020_o0,
			o0 => And249300_o0
		);
		Or249320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249300_o0,
			i1 => And249280_o0,
			o0 => Or249320_o0
		);
		And249340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249320_o0,
			i1 => Or210400_o0,
			o0 => And249340_o0
		);
		Or249360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i18,
			o0 => Or249360_o0
		);
		Or249380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or249360_o0,
			i1 => Not1040_o0,
			o0 => Or249380_o0
		);
		And249400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249380_o0,
			i1 => Xor2960_o0,
			o0 => And249400_o0
		);
		Or249420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210020_o0,
			i1 => i38,
			o0 => Or249420_o0
		);
		And249440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210420_o0,
			i1 => Nor21220_o0,
			o0 => And249440_o0
		);
		And249460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And249440_o0,
			i1 => Or249420_o0,
			o0 => And249460_o0
		);
		And249480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214120_o0,
			i1 => Not1280_o0,
			o0 => And249480_o0
		);
		Or249500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249480_o0,
			i1 => And215820_o0,
			o0 => Or249500_o0
		);
		Or249520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or249500_o0,
			i1 => And249460_o0,
			o0 => Or249520_o0
		);
		Or249540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or249520_o0,
			i1 => And249400_o0,
			o0 => Or249540_o0
		);
		Or249560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or249540_o0,
			i1 => i13,
			o0 => Or249560_o0
		);
		And249580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249560_o0,
			i1 => i12,
			o0 => And249580_o0
		);
		Or249600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21060_o0,
			i1 => Not2080_o0,
			o0 => Or249600_o0
		);
		And249620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249600_o0,
			i1 => Not28160_o0,
			o0 => And249620_o0
		);
		And249640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or219240_o0,
			i1 => Xor216140_o0,
			o0 => And249640_o0
		);
		Or249660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249640_o0,
			i1 => And23440_o0,
			o0 => Or249660_o0
		);
		Or249680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or249660_o0,
			i1 => And249620_o0,
			o0 => Or249680_o0
		);
		And249700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249680_o0,
			i1 => Not180_o0,
			o0 => And249700_o0
		);
		Or249720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249700_o0,
			i1 => And249580_o0,
			o0 => Or249720_o0
		);
		And249740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249720_o0,
			i1 => Not620_o0,
			o0 => And249740_o0
		);
		Or249760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or219240_o0,
			i1 => Not1040_o0,
			o0 => Or249760_o0
		);
		And249780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249760_o0,
			i1 => i18,
			o0 => And249780_o0
		);
		Or249800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249780_o0,
			i1 => And219340_o0,
			o0 => Or249800_o0
		);
		And249820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249800_o0,
			i1 => Not180_o0,
			o0 => And249820_o0
		);
		Or249840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And25700_o0,
			i1 => i12,
			o0 => Or249840_o0
		);
		And249860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249840_o0,
			i1 => i13,
			o0 => And249860_o0
		);
		And249880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Not1040_o0,
			o0 => And249880_o0
		);
		And249900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And249880_o0,
			i1 => Nand217420_o0,
			o0 => And249900_o0
		);
		Or249920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249900_o0,
			i1 => And249860_o0,
			o0 => Or249920_o0
		);
		And249940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or249920_o0,
			i1 => Not1280_o0,
			o0 => And249940_o0
		);
		And249960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or228180_o0,
			i1 => And23080_o0,
			o0 => And249960_o0
		);
		And249980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22480_o0,
			i1 => i12,
			o0 => And249980_o0
		);
		Or250000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And249980_o0,
			i1 => And249960_o0,
			o0 => Or250000_o0
		);
		Or250020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250000_o0,
			i1 => And249940_o0,
			o0 => Or250020_o0
		);
		Or250040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250020_o0,
			i1 => And249820_o0,
			o0 => Or250040_o0
		);
		And250060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250040_o0,
			i1 => i15,
			o0 => And250060_o0
		);
		Or250080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250060_o0,
			i1 => And249740_o0,
			o0 => Or250080_o0
		);
		And250100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250080_o0,
			i1 => Not540_o0,
			o0 => And250100_o0
		);
		And250120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => And2240_o0,
			o0 => And250120_o0
		);
		Or250140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250120_o0,
			i1 => i16,
			o0 => Or250140_o0
		);
		And250160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211940_o0,
			i1 => And211020_o0,
			o0 => And250160_o0
		);
		And250180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And250160_o0,
			i1 => Or250140_o0,
			o0 => And250180_o0
		);
		Or250200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250180_o0,
			i1 => And250100_o0,
			o0 => Or250200_o0
		);
		And250220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250200_o0,
			i1 => i40,
			o0 => And250220_o0
		);
		Or250240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250220_o0,
			i1 => And249340_o0,
			o0 => Or250240_o0
		);
		And250260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250240_o0,
			i1 => Not80_o0,
			o0 => And250260_o0
		);
		And250280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And244400_o0,
			i1 => i5,
			o0 => And250280_o0
		);
		And250300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor245680_o0,
			i1 => Not540_o0,
			o0 => And250300_o0
		);
		Nor250320 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor246000_o0,
			i1 => i5,
			o0 => Nor250320_o0
		);
		And250340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28120_o0,
			i1 => i5,
			o0 => And250340_o0
		);
		And250360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And250340_o0,
			i1 => And227280_o0,
			o0 => And250360_o0
		);
		Or250380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250360_o0,
			i1 => Nor250320_o0,
			o0 => Or250380_o0
		);
		Or250400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250380_o0,
			i1 => And250300_o0,
			o0 => Or250400_o0
		);
		And250420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225320_o0,
			i1 => i12,
			o0 => And250420_o0
		);
		Or250440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250420_o0,
			i1 => And239320_o0,
			o0 => Or250440_o0
		);
		And250460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i5,
			o0 => And250460_o0
		);
		And250480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And250460_o0,
			i1 => Or250440_o0,
			o0 => And250480_o0
		);
		And250500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And211940_o0,
			i1 => And24280_o0,
			o0 => And250500_o0
		);
		Or250520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250500_o0,
			i1 => And239880_o0,
			o0 => Or250520_o0
		);
		Or250540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250520_o0,
			i1 => And250480_o0,
			o0 => Or250540_o0
		);
		Or250560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250540_o0,
			i1 => Or250400_o0,
			o0 => Or250560_o0
		);
		Or250580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250560_o0,
			i1 => And250280_o0,
			o0 => Or250580_o0
		);
		And250600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250580_o0,
			i1 => And24040_o0,
			o0 => And250600_o0
		);
		Or250620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250600_o0,
			i1 => Nor233300_o0,
			o0 => Or250620_o0
		);
		Or250640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250620_o0,
			i1 => And250260_o0,
			o0 => Or250640_o0
		);
		And250660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250640_o0,
			i1 => Not160_o0,
			o0 => And250660_o0
		);
		And250680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247540_o0,
			i1 => i4,
			o0 => And250680_o0
		);
		Or250700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250680_o0,
			i1 => And250660_o0,
			o0 => Or250700_o0
		);
		And250720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250700_o0,
			i1 => Not140_o0,
			o0 => And250720_o0
		);
		And250740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248140_o0,
			i1 => i3,
			o0 => And250740_o0
		);
		Or250760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250740_o0,
			i1 => And250720_o0,
			o0 => Or250760_o0
		);
		And250780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250760_o0,
			i1 => Not120_o0,
			o0 => And250780_o0
		);
		And250800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248400_o0,
			i1 => i2,
			o0 => And250800_o0
		);
		Or250820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250800_o0,
			i1 => And250780_o0,
			o0 => Or250820_o0
		);
		And250840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250820_o0,
			i1 => Not100_o0,
			o0 => And250840_o0
		);
		Or250860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250840_o0,
			i1 => And230880_o0,
			o0 => Or250860_o0
		);
		And250880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250860_o0,
			i1 => Not60_o0,
			o0 => And250880_o0
		);
		And250900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248640_o0,
			i1 => And242020_o0,
			o0 => And250900_o0
		);
		Or250920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And250900_o0,
			i1 => And250880_o0,
			o0 => Or250920_o0
		);
		Or250940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250920_o0,
			i1 => i36,
			o0 => Or250940_o0
		);
		Or250960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250940_o0,
			i1 => i10,
			o0 => Or250960_o0
		);
		Or250980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or250960_o0,
			i1 => i9,
			o0 => Or250980_o0
		);
		And251000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or250980_o0,
			i1 => Not24960_o0,
			o0 => And251000_o0
		);
		Or251020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251000_o0,
			i1 => And235000_o0,
			o0 => Or251020_o0
		);
		And251040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251020_o0,
			i1 => Not12100_o0,
			o0 => And251040_o0
		);
		Or251060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251040_o0,
			i1 => And235080_o0,
			o0 => Or251060_o0
		);
		And251080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor26660_o0,
			i1 => Nor24920_o0,
			o0 => And251080_o0
		);
		And251100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => And23080_o0,
			o0 => And251100_o0
		);
		And251120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And251100_o0,
			i1 => And251080_o0,
			o0 => And251120_o0
		);
		And251140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And251120_o0,
			i1 => And23340_o0,
			o0 => And251140_o0
		);
		And251160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And251140_o0,
			i1 => And213280_o0,
			o0 => And251160_o0
		);
		And251180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And251140_o0,
			i1 => And23640_o0,
			o0 => And251180_o0
		);
		Or251200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251180_o0,
			i1 => i10,
			o0 => Or251200_o0
		);
		And251220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251200_o0,
			i1 => Nor23280_o0,
			o0 => And251220_o0
		);
		Or251240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And226340_o0,
			i1 => i13,
			o0 => Or251240_o0
		);
		And251260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251240_o0,
			i1 => i12,
			o0 => And251260_o0
		);
		Or251280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or228180_o0,
			i1 => And212900_o0,
			o0 => Or251280_o0
		);
		And251300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251280_o0,
			i1 => And23080_o0,
			o0 => And251300_o0
		);
		Or251320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251300_o0,
			i1 => Not180_o0,
			o0 => Or251320_o0
		);
		Or251340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or251320_o0,
			i1 => And251260_o0,
			o0 => Or251340_o0
		);
		And251360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251340_o0,
			i1 => i15,
			o0 => And251360_o0
		);
		Or251380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251360_o0,
			i1 => And245540_o0,
			o0 => Or251380_o0
		);
		And251400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251380_o0,
			i1 => Not80_o0,
			o0 => And251400_o0
		);
		Or251420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251400_o0,
			i1 => And246060_o0,
			o0 => Or251420_o0
		);
		Or251440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or251420_o0,
			i1 => Not24560_o0,
			o0 => Or251440_o0
		);
		And251460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251440_o0,
			i1 => Nor214960_o0,
			o0 => And251460_o0
		);
		Or251480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251460_o0,
			i1 => i8,
			o0 => Or251480_o0
		);
		And251500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251480_o0,
			i1 => Not540_o0,
			o0 => And251500_o0
		);
		Or251520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251500_o0,
			i1 => And247240_o0,
			o0 => Or251520_o0
		);
		And251540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251520_o0,
			i1 => Not160_o0,
			o0 => And251540_o0
		);
		Or251560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251540_o0,
			i1 => And247600_o0,
			o0 => Or251560_o0
		);
		And251580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251560_o0,
			i1 => Not140_o0,
			o0 => And251580_o0
		);
		Or251600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251580_o0,
			i1 => And248200_o0,
			o0 => Or251600_o0
		);
		And251620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251600_o0,
			i1 => Not120_o0,
			o0 => And251620_o0
		);
		Or251640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251620_o0,
			i1 => And248460_o0,
			o0 => Or251640_o0
		);
		And251660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251640_o0,
			i1 => Not100_o0,
			o0 => And251660_o0
		);
		Or251680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251660_o0,
			i1 => And248560_o0,
			o0 => Or251680_o0
		);
		And251700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251680_o0,
			i1 => Not60_o0,
			o0 => And251700_o0
		);
		Or251720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251700_o0,
			i1 => And248720_o0,
			o0 => Or251720_o0
		);
		And251740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251720_o0,
			i1 => Not3300_o0,
			o0 => And251740_o0
		);
		Or251760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251740_o0,
			i1 => And248800_o0,
			o0 => Or251760_o0
		);
		And251780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251760_o0,
			i1 => Not24960_o0,
			o0 => And251780_o0
		);
		Or251800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251780_o0,
			i1 => And248860_o0,
			o0 => Or251800_o0
		);
		And251820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251800_o0,
			i1 => Not20520_o0,
			o0 => And251820_o0
		);
		Or251840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251820_o0,
			i1 => And248940_o0,
			o0 => Or251840_o0
		);
		Xor251860 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => i9,
			o0 => Xor251860_o0
		);
		Or251880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Xor251860_o0,
			i1 => And220460_o0,
			o0 => Or251880_o0
		);
		And251900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or251880_o0,
			i1 => Not12100_o0,
			o0 => And251900_o0
		);
		And251920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220180_o0,
			i1 => i15,
			o0 => And251920_o0
		);
		And251940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2240_o0,
			i1 => Not620_o0,
			o0 => And251940_o0
		);
		Or251960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And251940_o0,
			i1 => And251920_o0,
			o0 => Or251960_o0
		);
		And251980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28040_o0,
			i1 => Nor21260_o0,
			o0 => And251980_o0
		);
		And252000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And251980_o0,
			i1 => And28160_o0,
			o0 => And252000_o0
		);
		Nor252020 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i14,
			o0 => Nor252020_o0
		);
		And252040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor252020_o0,
			i1 => And23080_o0,
			o0 => And252040_o0
		);
		And252060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252040_o0,
			i1 => And23340_o0,
			o0 => And252060_o0
		);
		And252080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252060_o0,
			i1 => And252000_o0,
			o0 => And252080_o0
		);
		And252100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252080_o0,
			i1 => Or251960_o0,
			o0 => And252100_o0
		);
		Or252120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252100_o0,
			i1 => i10,
			o0 => Or252120_o0
		);
		And252140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252120_o0,
			i1 => Not20520_o0,
			o0 => And252140_o0
		);
		Or252160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252140_o0,
			i1 => And212160_o0,
			o0 => Or252160_o0
		);
		And252180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252160_o0,
			i1 => Not12100_o0,
			o0 => And252180_o0
		);
		Or252200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nand223780_o0,
			i1 => Not1080_o0,
			o0 => Or252200_o0
		);
		And252220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252200_o0,
			i1 => And23020_o0,
			o0 => And252220_o0
		);
		Or252240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252220_o0,
			i1 => And245840_o0,
			o0 => Or252240_o0
		);
		And252260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252240_o0,
			i1 => Nor22900_o0,
			o0 => And252260_o0
		);
		Or252280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252260_o0,
			i1 => Or245780_o0,
			o0 => Or252280_o0
		);
		Or252300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or252280_o0,
			i1 => And251260_o0,
			o0 => Or252300_o0
		);
		And252320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252300_o0,
			i1 => i15,
			o0 => And252320_o0
		);
		Or252340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252320_o0,
			i1 => And245540_o0,
			o0 => Or252340_o0
		);
		And252360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252340_o0,
			i1 => Not80_o0,
			o0 => And252360_o0
		);
		Or252380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252360_o0,
			i1 => And246060_o0,
			o0 => Or252380_o0
		);
		Or252400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or252380_o0,
			i1 => Not24560_o0,
			o0 => Or252400_o0
		);
		And252420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214960_o0,
			i1 => Not24960_o0,
			o0 => And252420_o0
		);
		And252440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252420_o0,
			i1 => Or252400_o0,
			o0 => And252440_o0
		);
		Or252460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252440_o0,
			i1 => i8,
			o0 => Or252460_o0
		);
		And252480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252460_o0,
			i1 => Not540_o0,
			o0 => And252480_o0
		);
		And252500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227400_o0,
			i1 => Nor23320_o0,
			o0 => And252500_o0
		);
		And252520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252500_o0,
			i1 => Or247200_o0,
			o0 => And252520_o0
		);
		Or252540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252520_o0,
			i1 => And252480_o0,
			o0 => Or252540_o0
		);
		And252560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252540_o0,
			i1 => Not160_o0,
			o0 => And252560_o0
		);
		And252580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And247560_o0,
			i1 => Nor23320_o0,
			o0 => And252580_o0
		);
		And252600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252580_o0,
			i1 => And247540_o0,
			o0 => And252600_o0
		);
		Or252620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252600_o0,
			i1 => And252560_o0,
			o0 => Or252620_o0
		);
		And252640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252620_o0,
			i1 => Not140_o0,
			o0 => And252640_o0
		);
		And252660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248160_o0,
			i1 => Nor23320_o0,
			o0 => And252660_o0
		);
		And252680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252660_o0,
			i1 => And248140_o0,
			o0 => And252680_o0
		);
		Or252700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252680_o0,
			i1 => And252640_o0,
			o0 => Or252700_o0
		);
		And252720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252700_o0,
			i1 => Not120_o0,
			o0 => And252720_o0
		);
		And252740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248420_o0,
			i1 => Nor23320_o0,
			o0 => And252740_o0
		);
		And252760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252740_o0,
			i1 => And248400_o0,
			o0 => And252760_o0
		);
		Or252780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252760_o0,
			i1 => And252720_o0,
			o0 => Or252780_o0
		);
		And252800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252780_o0,
			i1 => Not100_o0,
			o0 => And252800_o0
		);
		And252820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And248520_o0,
			i1 => Nor23320_o0,
			o0 => And252820_o0
		);
		And252840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252820_o0,
			i1 => And230860_o0,
			o0 => And252840_o0
		);
		Or252860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252840_o0,
			i1 => And252800_o0,
			o0 => Or252860_o0
		);
		And252880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252860_o0,
			i1 => Not60_o0,
			o0 => And252880_o0
		);
		And252900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor248660_o0,
			i1 => Nor23320_o0,
			o0 => And252900_o0
		);
		And252920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252900_o0,
			i1 => And23180_o0,
			o0 => And252920_o0
		);
		And252940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252920_o0,
			i1 => And248640_o0,
			o0 => And252940_o0
		);
		Or252960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And252940_o0,
			i1 => And252880_o0,
			o0 => Or252960_o0
		);
		And252980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or252960_o0,
			i1 => Not3300_o0,
			o0 => And252980_o0
		);
		And253000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => Not24960_o0,
			o0 => And253000_o0
		);
		And253020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And253000_o0,
			i1 => Nor214960_o0,
			o0 => And253020_o0
		);
		Or253040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253020_o0,
			i1 => And252980_o0,
			o0 => Or253040_o0
		);
		And253060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253040_o0,
			i1 => Not20520_o0,
			o0 => And253060_o0
		);
		Or253080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253060_o0,
			i1 => And248940_o0,
			o0 => Or253080_o0
		);
		And253100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244960_o0,
			i1 => i17,
			o0 => And253100_o0
		);
		Or253120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not1080_o0,
			i1 => i16,
			o0 => Or253120_o0
		);
		And253140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253120_o0,
			i1 => Not1040_o0,
			o0 => And253140_o0
		);
		Or253160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253140_o0,
			i1 => And253100_o0,
			o0 => Or253160_o0
		);
		And253180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253160_o0,
			i1 => Not2080_o0,
			o0 => And253180_o0
		);
		Or253200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253180_o0,
			i1 => Or245420_o0,
			o0 => Or253200_o0
		);
		And253220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253200_o0,
			i1 => i12,
			o0 => And253220_o0
		);
		Or253240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253220_o0,
			i1 => And245500_o0,
			o0 => Or253240_o0
		);
		And253260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253240_o0,
			i1 => Not620_o0,
			o0 => And253260_o0
		);
		And253280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215260_o0,
			i1 => Not1040_o0,
			o0 => And253280_o0
		);
		And253300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And253280_o0,
			i1 => And232100_o0,
			o0 => And253300_o0
		);
		Or253320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253300_o0,
			i1 => i13,
			o0 => Or253320_o0
		);
		And253340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253320_o0,
			i1 => i12,
			o0 => And253340_o0
		);
		Or253360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253340_o0,
			i1 => Or252280_o0,
			o0 => Or253360_o0
		);
		And253380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253360_o0,
			i1 => i15,
			o0 => And253380_o0
		);
		Or253400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253380_o0,
			i1 => And253260_o0,
			o0 => Or253400_o0
		);
		And253420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253400_o0,
			i1 => Not80_o0,
			o0 => And253420_o0
		);
		Or253440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253420_o0,
			i1 => And246060_o0,
			o0 => Or253440_o0
		);
		Or253460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or253440_o0,
			i1 => Not24560_o0,
			o0 => Or253460_o0
		);
		And253480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253460_o0,
			i1 => And252420_o0,
			o0 => And253480_o0
		);
		Or253500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253480_o0,
			i1 => i8,
			o0 => Or253500_o0
		);
		And253520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253500_o0,
			i1 => Not540_o0,
			o0 => And253520_o0
		);
		Or253540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253520_o0,
			i1 => And252520_o0,
			o0 => Or253540_o0
		);
		And253560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253540_o0,
			i1 => Not160_o0,
			o0 => And253560_o0
		);
		Or253580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253560_o0,
			i1 => And252600_o0,
			o0 => Or253580_o0
		);
		And253600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253580_o0,
			i1 => Not140_o0,
			o0 => And253600_o0
		);
		Or253620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253600_o0,
			i1 => And252680_o0,
			o0 => Or253620_o0
		);
		And253640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253620_o0,
			i1 => Not120_o0,
			o0 => And253640_o0
		);
		Or253660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253640_o0,
			i1 => And252760_o0,
			o0 => Or253660_o0
		);
		And253680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253660_o0,
			i1 => Not100_o0,
			o0 => And253680_o0
		);
		Or253700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253680_o0,
			i1 => And252840_o0,
			o0 => Or253700_o0
		);
		And253720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253700_o0,
			i1 => Not60_o0,
			o0 => And253720_o0
		);
		Or253740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253720_o0,
			i1 => And252940_o0,
			o0 => Or253740_o0
		);
		And253760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253740_o0,
			i1 => Not3300_o0,
			o0 => And253760_o0
		);
		Or253780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253760_o0,
			i1 => And253020_o0,
			o0 => Or253780_o0
		);
		And253800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253780_o0,
			i1 => Not20520_o0,
			o0 => And253800_o0
		);
		Or253820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253800_o0,
			i1 => And248940_o0,
			o0 => Or253820_o0
		);
		And253840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor212260_o0,
			i1 => And25420_o0,
			o0 => And253840_o0
		);
		And253860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => Not620_o0,
			o0 => And253860_o0
		);
		Or253880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253860_o0,
			i1 => And253840_o0,
			o0 => Or253880_o0
		);
		And253900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or253880_o0,
			i1 => Not1500_o0,
			o0 => And253900_o0
		);
		Or253920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And253900_o0,
			i1 => And251940_o0,
			o0 => Or253920_o0
		);
		And253940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23280_o0,
			i1 => Nor21140_o0,
			o0 => And253940_o0
		);
		And253960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And253940_o0,
			i1 => Nor23600_o0,
			o0 => And253960_o0
		);
		And253980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And252040_o0,
			i1 => And251980_o0,
			o0 => And253980_o0
		);
		And254000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And253980_o0,
			i1 => And23340_o0,
			o0 => And254000_o0
		);
		And254020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254000_o0,
			i1 => And253960_o0,
			o0 => And254020_o0
		);
		And254040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254020_o0,
			i1 => Or253920_o0,
			o0 => And254040_o0
		);
		And254060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218540_o0,
			i1 => i0,
			o0 => And254060_o0
		);
		Or254080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => Not1040_o0,
			o0 => Or254080_o0
		);
		And254100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254080_o0,
			i1 => Not1080_o0,
			o0 => And254100_o0
		);
		Or254120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254100_o0,
			i1 => And215080_o0,
			o0 => Or254120_o0
		);
		And254140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor237580_o0,
			i1 => And223380_o0,
			o0 => And254140_o0
		);
		And254160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254140_o0,
			i1 => Or254120_o0,
			o0 => And254160_o0
		);
		Or254180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254160_o0,
			i1 => And254060_o0,
			o0 => Or254180_o0
		);
		And254200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254180_o0,
			i1 => i16,
			o0 => And254200_o0
		);
		And254220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1500_o0,
			i1 => i3,
			o0 => And254220_o0
		);
		And254240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i18,
			i1 => Not140_o0,
			o0 => And254240_o0
		);
		And254260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254240_o0,
			i1 => And224580_o0,
			o0 => And254260_o0
		);
		Or254280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254260_o0,
			i1 => And254220_o0,
			o0 => Or254280_o0
		);
		And254300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i15,
			i1 => Not60_o0,
			o0 => And254300_o0
		);
		And254320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254300_o0,
			i1 => And21940_o0,
			o0 => And254320_o0
		);
		And254340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254320_o0,
			i1 => Or254280_o0,
			o0 => And254340_o0
		);
		Or254360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254340_o0,
			i1 => And254200_o0,
			o0 => Or254360_o0
		);
		And254380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254360_o0,
			i1 => Not180_o0,
			o0 => And254380_o0
		);
		And254400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i26,
			i1 => i25,
			o0 => And254400_o0
		);
		And254420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254400_o0,
			i1 => And25740_o0,
			o0 => And254420_o0
		);
		Or254440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254420_o0,
			i1 => i15,
			o0 => Or254440_o0
		);
		And254460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25840_o0,
			i1 => i28,
			o0 => And254460_o0
		);
		And254480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254460_o0,
			i1 => Nor237580_o0,
			o0 => And254480_o0
		);
		And254500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254480_o0,
			i1 => Or254440_o0,
			o0 => And254500_o0
		);
		Or254520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254500_o0,
			i1 => And254380_o0,
			o0 => Or254520_o0
		);
		And254540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254520_o0,
			i1 => i13,
			o0 => And254540_o0
		);
		And254560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor216140_o0,
			i1 => Xor2200_o0,
			o0 => And254560_o0
		);
		And254580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254560_o0,
			i1 => And26520_o0,
			o0 => And254580_o0
		);
		And254600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29740_o0,
			i1 => And26680_o0,
			o0 => And254600_o0
		);
		And254620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => Not1280_o0,
			o0 => And254620_o0
		);
		And254640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254620_o0,
			i1 => And245220_o0,
			o0 => And254640_o0
		);
		And254660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254640_o0,
			i1 => And254600_o0,
			o0 => And254660_o0
		);
		Or254680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254660_o0,
			i1 => And254580_o0,
			o0 => Or254680_o0
		);
		And254700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => Not60_o0,
			o0 => And254700_o0
		);
		And254720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => Not2080_o0,
			o0 => And254720_o0
		);
		And254740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254720_o0,
			i1 => And254700_o0,
			o0 => And254740_o0
		);
		And254760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254740_o0,
			i1 => Or254680_o0,
			o0 => And254760_o0
		);
		Or254780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254760_o0,
			i1 => And254540_o0,
			o0 => Or254780_o0
		);
		And254800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254780_o0,
			i1 => Not540_o0,
			o0 => And254800_o0
		);
		And254820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => i23,
			o0 => And254820_o0
		);
		Nor254840 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Not9580_o0,
			i1 => i26,
			o0 => Nor254840_o0
		);
		And254860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor254840_o0,
			i1 => And254820_o0,
			o0 => And254860_o0
		);
		Or254880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254860_o0,
			i1 => Nor218040_o0,
			o0 => Or254880_o0
		);
		And254900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254880_o0,
			i1 => i22,
			o0 => And254900_o0
		);
		Or254920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254900_o0,
			i1 => And218160_o0,
			o0 => Or254920_o0
		);
		And254940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or254920_o0,
			i1 => And29560_o0,
			o0 => And254940_o0
		);
		Or254960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And254940_o0,
			i1 => And218280_o0,
			o0 => Or254960_o0
		);
		And254980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => And21940_o0,
			o0 => And254980_o0
		);
		And255000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240360_o0,
			i1 => Nor211040_o0,
			o0 => And255000_o0
		);
		And255020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255000_o0,
			i1 => And254700_o0,
			o0 => And255020_o0
		);
		And255040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255020_o0,
			i1 => And254980_o0,
			o0 => And255040_o0
		);
		And255060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255040_o0,
			i1 => Or254960_o0,
			o0 => And255060_o0
		);
		Or255080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255060_o0,
			i1 => And254800_o0,
			o0 => Or255080_o0
		);
		And255100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255080_o0,
			i1 => Not80_o0,
			o0 => And255100_o0
		);
		And255120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28060_o0,
			i1 => i16,
			o0 => And255120_o0
		);
		And255140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255120_o0,
			i1 => And28040_o0,
			o0 => And255140_o0
		);
		And255160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237600_o0,
			i1 => And222800_o0,
			o0 => And255160_o0
		);
		And255180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255160_o0,
			i1 => And255140_o0,
			o0 => And255180_o0
		);
		Or255200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255180_o0,
			i1 => And255100_o0,
			o0 => Or255200_o0
		);
		And255220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255200_o0,
			i1 => Not120_o0,
			o0 => And255220_o0
		);
		And255240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor237580_o0,
			i1 => i2,
			o0 => And255240_o0
		);
		And255260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255240_o0,
			i1 => And219040_o0,
			o0 => And255260_o0
		);
		Or255280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255260_o0,
			i1 => And255220_o0,
			o0 => Or255280_o0
		);
		And255300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255280_o0,
			i1 => Not160_o0,
			o0 => And255300_o0
		);
		And255320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218560_o0,
			i1 => And29940_o0,
			o0 => And255320_o0
		);
		And255340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26680_o0,
			i1 => i17,
			o0 => And255340_o0
		);
		And255360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255340_o0,
			i1 => Nor229280_o0,
			o0 => And255360_o0
		);
		And255380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255360_o0,
			i1 => And234580_o0,
			o0 => And255380_o0
		);
		Or255400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255380_o0,
			i1 => And255320_o0,
			o0 => Or255400_o0
		);
		And255420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215260_o0,
			i1 => i18,
			o0 => And255420_o0
		);
		And255440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24560_o0,
			i1 => Nor23200_o0,
			o0 => And255440_o0
		);
		And255460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255440_o0,
			i1 => And254700_o0,
			o0 => And255460_o0
		);
		And255480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255460_o0,
			i1 => And255420_o0,
			o0 => And255480_o0
		);
		And255500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255480_o0,
			i1 => Or255400_o0,
			o0 => And255500_o0
		);
		Or255520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255500_o0,
			i1 => And255300_o0,
			o0 => Or255520_o0
		);
		Nor255540 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			i1 => i8,
			o0 => Nor255540_o0
		);
		And255560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor255540_o0,
			i1 => Nor212700_o0,
			o0 => And255560_o0
		);
		And255580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255560_o0,
			i1 => Nor234860_o0,
			o0 => And255580_o0
		);
		And255600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255580_o0,
			i1 => Or255520_o0,
			o0 => And255600_o0
		);
		And255620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219060_o0,
			i1 => Not540_o0,
			o0 => And255620_o0
		);
		And255640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255620_o0,
			i1 => And221440_o0,
			o0 => And255640_o0
		);
		And255660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233760_o0,
			i1 => Not9580_o0,
			o0 => And255660_o0
		);
		And255680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255660_o0,
			i1 => And243960_o0,
			o0 => And255680_o0
		);
		Or255700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255680_o0,
			i1 => And255640_o0,
			o0 => Or255700_o0
		);
		And255720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255700_o0,
			i1 => Not7120_o0,
			o0 => And255720_o0
		);
		And255740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And244800_o0,
			i1 => And233760_o0,
			o0 => And255740_o0
		);
		And255760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255740_o0,
			i1 => And243960_o0,
			o0 => And255760_o0
		);
		Or255780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255760_o0,
			i1 => And255720_o0,
			o0 => Or255780_o0
		);
		And255800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255780_o0,
			i1 => And29560_o0,
			o0 => And255800_o0
		);
		And255820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24400_o0,
			i1 => i2,
			o0 => And255820_o0
		);
		And255840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255820_o0,
			i1 => And230320_o0,
			o0 => And255840_o0
		);
		Or255860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255840_o0,
			i1 => And255800_o0,
			o0 => Or255860_o0
		);
		And255880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255860_o0,
			i1 => Not620_o0,
			o0 => And255880_o0
		);
		And255900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246320_o0,
			i1 => Not540_o0,
			o0 => And255900_o0
		);
		And255920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255900_o0,
			i1 => Nor21140_o0,
			o0 => And255920_o0
		);
		Or255940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And255920_o0,
			i1 => And255880_o0,
			o0 => Or255940_o0
		);
		And255960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or255940_o0,
			i1 => And215060_o0,
			o0 => And255960_o0
		);
		And255980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => And25420_o0,
			o0 => And255980_o0
		);
		And256000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255980_o0,
			i1 => And242460_o0,
			o0 => And256000_o0
		);
		Or256020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256000_o0,
			i1 => And255960_o0,
			o0 => Or256020_o0
		);
		And256040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256020_o0,
			i1 => i17,
			o0 => And256040_o0
		);
		And256060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22940_o0,
			i1 => Nor21140_o0,
			o0 => And256060_o0
		);
		And256080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222120_o0,
			i1 => And212880_o0,
			o0 => And256080_o0
		);
		And256100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256080_o0,
			i1 => And256060_o0,
			o0 => And256100_o0
		);
		Or256120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256100_o0,
			i1 => And256040_o0,
			o0 => Or256120_o0
		);
		And256140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256120_o0,
			i1 => Not1280_o0,
			o0 => And256140_o0
		);
		And256160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21980_o0,
			i1 => Nor21140_o0,
			o0 => And256160_o0
		);
		And256180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256160_o0,
			i1 => And210420_o0,
			o0 => And256180_o0
		);
		And256200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256180_o0,
			i1 => And224600_o0,
			o0 => And256200_o0
		);
		Or256220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256200_o0,
			i1 => And256140_o0,
			o0 => Or256220_o0
		);
		And256240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256220_o0,
			i1 => Not2080_o0,
			o0 => And256240_o0
		);
		And256260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i34,
			i1 => i33,
			o0 => And256260_o0
		);
		And256280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256260_o0,
			i1 => i13,
			o0 => And256280_o0
		);
		And256300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29420_o0,
			i1 => And2560_o0,
			o0 => And256300_o0
		);
		And256320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256300_o0,
			i1 => Nor21140_o0,
			o0 => And256320_o0
		);
		And256340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256320_o0,
			i1 => And256280_o0,
			o0 => And256340_o0
		);
		Or256360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256340_o0,
			i1 => And256240_o0,
			o0 => Or256360_o0
		);
		And256380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256360_o0,
			i1 => Not80_o0,
			o0 => And256380_o0
		);
		And256400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246320_o0,
			i1 => And223260_o0,
			o0 => And256400_o0
		);
		And256420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256400_o0,
			i1 => And242460_o0,
			o0 => And256420_o0
		);
		Or256440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256420_o0,
			i1 => And256380_o0,
			o0 => Or256440_o0
		);
		And256460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256440_o0,
			i1 => i12,
			o0 => And256460_o0
		);
		And256480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => Nor21140_o0,
			o0 => And256480_o0
		);
		And256500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246320_o0,
			i1 => Nor232220_o0,
			o0 => And256500_o0
		);
		And256520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256500_o0,
			i1 => And256480_o0,
			o0 => And256520_o0
		);
		Or256540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256520_o0,
			i1 => And256460_o0,
			o0 => Or256540_o0
		);
		And256560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256540_o0,
			i1 => Not160_o0,
			o0 => And256560_o0
		);
		And256580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24560_o0,
			i1 => And26040_o0,
			o0 => And256580_o0
		);
		And256600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256580_o0,
			i1 => And234620_o0,
			o0 => And256600_o0
		);
		And256620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256600_o0,
			i1 => And234600_o0,
			o0 => And256620_o0
		);
		Or256640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256620_o0,
			i1 => And256560_o0,
			o0 => Or256640_o0
		);
		And256660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23600_o0,
			i1 => Nor23280_o0,
			o0 => And256660_o0
		);
		And256680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256660_o0,
			i1 => And23340_o0,
			o0 => And256680_o0
		);
		And256700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256680_o0,
			i1 => Or256640_o0,
			o0 => And256700_o0
		);
		And256720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i26,
			o0 => And256720_o0
		);
		And256740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9580_o0,
			i1 => i25,
			o0 => And256740_o0
		);
		Or256760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256740_o0,
			i1 => And256720_o0,
			o0 => Or256760_o0
		);
		And256780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256760_o0,
			i1 => And254820_o0,
			o0 => And256780_o0
		);
		And256800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9540_o0,
			i1 => i12,
			o0 => And256800_o0
		);
		And256820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256800_o0,
			i1 => And234540_o0,
			o0 => And256820_o0
		);
		And256840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256820_o0,
			i1 => And229420_o0,
			o0 => And256840_o0
		);
		And256860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256840_o0,
			i1 => And256780_o0,
			o0 => And256860_o0
		);
		Nor256880 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i3,
			o0 => Nor256880_o0
		);
		And256900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor256880_o0,
			i1 => And24040_o0,
			o0 => And256900_o0
		);
		Or256920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256900_o0,
			i1 => And256860_o0,
			o0 => Or256920_o0
		);
		And256940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or256920_o0,
			i1 => Not1500_o0,
			o0 => And256940_o0
		);
		And256960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => i14,
			o0 => And256960_o0
		);
		And256980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256960_o0,
			i1 => Nor256880_o0,
			o0 => And256980_o0
		);
		Or257000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And256980_o0,
			i1 => And256940_o0,
			o0 => Or257000_o0
		);
		And257020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257000_o0,
			i1 => Not620_o0,
			o0 => And257020_o0
		);
		And257040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246340_o0,
			i1 => Not140_o0,
			o0 => And257040_o0
		);
		Or257060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257040_o0,
			i1 => And257020_o0,
			o0 => Or257060_o0
		);
		And257080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257060_o0,
			i1 => Not1280_o0,
			o0 => And257080_o0
		);
		And257100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246440_o0,
			i1 => Not140_o0,
			o0 => And257100_o0
		);
		Or257120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257100_o0,
			i1 => And257080_o0,
			o0 => Or257120_o0
		);
		And257140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257120_o0,
			i1 => i18,
			o0 => And257140_o0
		);
		And257160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246520_o0,
			i1 => Not1080_o0,
			o0 => And257160_o0
		);
		And257180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257160_o0,
			i1 => Not140_o0,
			o0 => And257180_o0
		);
		Or257200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257180_o0,
			i1 => And257140_o0,
			o0 => Or257200_o0
		);
		And257220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257200_o0,
			i1 => i17,
			o0 => And257220_o0
		);
		Nor257240 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i3,
			o0 => Nor257240_o0
		);
		And257260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor257240_o0,
			i1 => And246640_o0,
			o0 => And257260_o0
		);
		Or257280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257260_o0,
			i1 => And257220_o0,
			o0 => Or257280_o0
		);
		And257300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257280_o0,
			i1 => Not2080_o0,
			o0 => And257300_o0
		);
		And257320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => i40,
			o0 => And257320_o0
		);
		And257340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257320_o0,
			i1 => And24140_o0,
			o0 => And257340_o0
		);
		And257360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257340_o0,
			i1 => Or233140_o0,
			o0 => And257360_o0
		);
		Or257380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257360_o0,
			i1 => And257300_o0,
			o0 => Or257380_o0
		);
		And257400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257380_o0,
			i1 => i5,
			o0 => And257400_o0
		);
		And257420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => Not1280_o0,
			o0 => And257420_o0
		);
		And257440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257420_o0,
			i1 => Xor216140_o0,
			o0 => And257440_o0
		);
		And257460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => i16,
			o0 => And257460_o0
		);
		And257480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257460_o0,
			i1 => And212560_o0,
			o0 => And257480_o0
		);
		Or257500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257480_o0,
			i1 => And257440_o0,
			o0 => Or257500_o0
		);
		And257520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257500_o0,
			i1 => i17,
			o0 => And257520_o0
		);
		Or257540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219800_o0,
			i1 => i14,
			o0 => Or257540_o0
		);
		And257560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257540_o0,
			i1 => Not2080_o0,
			o0 => And257560_o0
		);
		And257580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => i20,
			o0 => And257580_o0
		);
		And257600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And236820_o0,
			i1 => And234540_o0,
			o0 => And257600_o0
		);
		And257620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257600_o0,
			i1 => And257580_o0,
			o0 => And257620_o0
		);
		Or257640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257620_o0,
			i1 => And257560_o0,
			o0 => Or257640_o0
		);
		Or257660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or257640_o0,
			i1 => And257520_o0,
			o0 => Or257660_o0
		);
		And257680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257660_o0,
			i1 => i12,
			o0 => And257680_o0
		);
		And257700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244160_o0,
			i1 => i14,
			o0 => And257700_o0
		);
		And257720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21060_o0,
			i1 => And2240_o0,
			o0 => And257720_o0
		);
		Or257740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257720_o0,
			i1 => Not1280_o0,
			o0 => Or257740_o0
		);
		And257760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257740_o0,
			i1 => And23520_o0,
			o0 => And257760_o0
		);
		Or257780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257760_o0,
			i1 => And257700_o0,
			o0 => Or257780_o0
		);
		And257800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257780_o0,
			i1 => Not180_o0,
			o0 => And257800_o0
		);
		Or257820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257800_o0,
			i1 => And257680_o0,
			o0 => Or257820_o0
		);
		And257840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257820_o0,
			i1 => Not620_o0,
			o0 => And257840_o0
		);
		And257860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => And23080_o0,
			o0 => And257860_o0
		);
		And257880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257860_o0,
			i1 => And22920_o0,
			o0 => And257880_o0
		);
		Or257900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257880_o0,
			i1 => And257840_o0,
			o0 => Or257900_o0
		);
		And257920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or257900_o0,
			i1 => And26520_o0,
			o0 => And257920_o0
		);
		And257940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i3,
			o0 => And257940_o0
		);
		And257960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257940_o0,
			i1 => Nor29260_o0,
			o0 => And257960_o0
		);
		And257980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257960_o0,
			i1 => And23060_o0,
			o0 => And257980_o0
		);
		Or258000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And257980_o0,
			i1 => And257920_o0,
			o0 => Or258000_o0
		);
		And258020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258000_o0,
			i1 => Not540_o0,
			o0 => And258020_o0
		);
		Or258040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258020_o0,
			i1 => And257400_o0,
			o0 => Or258040_o0
		);
		And258060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258040_o0,
			i1 => Not60_o0,
			o0 => And258060_o0
		);
		And258080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26760_o0,
			i1 => And23100_o0,
			o0 => And258080_o0
		);
		And258100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And258080_o0,
			i1 => And214680_o0,
			o0 => And258100_o0
		);
		Or258120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258100_o0,
			i1 => And258060_o0,
			o0 => Or258120_o0
		);
		And258140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor220340_o0,
			i1 => Nor22060_o0,
			o0 => And258140_o0
		);
		And258160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And258140_o0,
			i1 => And215000_o0,
			o0 => And258160_o0
		);
		And258180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And258160_o0,
			i1 => Or258120_o0,
			o0 => And258180_o0
		);
		And258200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or29840_o0,
			i1 => Or25540_o0,
			o0 => And258200_o0
		);
		Or258220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233680_o0,
			i1 => Nand210560_o0,
			o0 => Or258220_o0
		);
		And258240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258220_o0,
			i1 => i27,
			o0 => And258240_o0
		);
		And258260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210560_o0,
			i1 => Nor29640_o0,
			o0 => And258260_o0
		);
		Or258280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258260_o0,
			i1 => And258240_o0,
			o0 => Or258280_o0
		);
		And258300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258280_o0,
			i1 => And26520_o0,
			o0 => And258300_o0
		);
		Or258320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258300_o0,
			i1 => And258200_o0,
			o0 => Or258320_o0
		);
		And258340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258320_o0,
			i1 => Not540_o0,
			o0 => And258340_o0
		);
		And258360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256780_o0,
			i1 => i3,
			o0 => And258360_o0
		);
		Nor258380 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i23,
			i1 => i3,
			o0 => Nor258380_o0
		);
		And258400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor258380_o0,
			i1 => And221240_o0,
			o0 => And258400_o0
		);
		Or258420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258400_o0,
			i1 => And258360_o0,
			o0 => Or258420_o0
		);
		And258440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258420_o0,
			i1 => i22,
			o0 => And258440_o0
		);
		And258460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217780_o0,
			i1 => i27,
			o0 => And258460_o0
		);
		And258480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And258460_o0,
			i1 => Nand210640_o0,
			o0 => And258480_o0
		);
		Nor258500 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			i1 => i3,
			o0 => Nor258500_o0
		);
		And258520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor258500_o0,
			i1 => And221240_o0,
			o0 => And258520_o0
		);
		Or258540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258520_o0,
			i1 => Nor247900_o0,
			o0 => Or258540_o0
		);
		Or258560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or258540_o0,
			i1 => And258480_o0,
			o0 => Or258560_o0
		);
		Or258580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or258560_o0,
			i1 => And258440_o0,
			o0 => Or258580_o0
		);
		And258600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258580_o0,
			i1 => i5,
			o0 => And258600_o0
		);
		Or258620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258600_o0,
			i1 => And258340_o0,
			o0 => Or258620_o0
		);
		And258640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258620_o0,
			i1 => Not160_o0,
			o0 => And258640_o0
		);
		And258660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i4,
			o0 => And258660_o0
		);
		Or258680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => Not140_o0,
			o0 => Or258680_o0
		);
		And258700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258680_o0,
			i1 => Nand210560_o0,
			o0 => And258700_o0
		);
		And258720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227520_o0,
			i1 => And217780_o0,
			o0 => And258720_o0
		);
		Or258740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258720_o0,
			i1 => And258700_o0,
			o0 => Or258740_o0
		);
		And258760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258740_o0,
			i1 => Not7120_o0,
			o0 => And258760_o0
		);
		And258780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227520_o0,
			i1 => And210740_o0,
			o0 => And258780_o0
		);
		Or258800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258780_o0,
			i1 => And258760_o0,
			o0 => Or258800_o0
		);
		And258820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258800_o0,
			i1 => And258660_o0,
			o0 => And258820_o0
		);
		Or258840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258820_o0,
			i1 => And258640_o0,
			o0 => Or258840_o0
		);
		And258860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258840_o0,
			i1 => Not9540_o0,
			o0 => And258860_o0
		);
		And258880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2560_o0,
			i1 => i20,
			o0 => And258880_o0
		);
		And258900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And258880_o0,
			i1 => Nor22600_o0,
			o0 => And258900_o0
		);
		Or258920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258900_o0,
			i1 => And258860_o0,
			o0 => Or258920_o0
		);
		And258940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258920_o0,
			i1 => i21,
			o0 => And258940_o0
		);
		And258960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or223040_o0,
			i1 => i27,
			o0 => And258960_o0
		);
		And258980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor217900_o0,
			i1 => Or210400_o0,
			o0 => And258980_o0
		);
		Or259000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And258980_o0,
			i1 => And258960_o0,
			o0 => Or259000_o0
		);
		And259020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259000_o0,
			i1 => Not140_o0,
			o0 => And259020_o0
		);
		And259040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9580_o0,
			i1 => i5,
			o0 => And259040_o0
		);
		And259060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259040_o0,
			i1 => And224200_o0,
			o0 => And259060_o0
		);
		Or259080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259060_o0,
			i1 => And259020_o0,
			o0 => Or259080_o0
		);
		And259100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259080_o0,
			i1 => And210540_o0,
			o0 => And259100_o0
		);
		Or259120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259100_o0,
			i1 => And258940_o0,
			o0 => Or259120_o0
		);
		And259140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259120_o0,
			i1 => Not120_o0,
			o0 => And259140_o0
		);
		Or259160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And218900_o0,
			i1 => And210540_o0,
			o0 => Or259160_o0
		);
		And259180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259160_o0,
			i1 => i27,
			o0 => And259180_o0
		);
		And259200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259180_o0,
			i1 => And219080_o0,
			o0 => And259200_o0
		);
		Or259220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259200_o0,
			i1 => And259140_o0,
			o0 => Or259220_o0
		);
		And259240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => And23080_o0,
			o0 => And259240_o0
		);
		And259260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259240_o0,
			i1 => And218980_o0,
			o0 => And259260_o0
		);
		And259280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259260_o0,
			i1 => And256680_o0,
			o0 => And259280_o0
		);
		And259300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259280_o0,
			i1 => Or259220_o0,
			o0 => And259300_o0
		);
		Or259320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And216540_o0,
			i1 => Or210620_o0,
			o0 => Or259320_o0
		);
		Or259340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or259320_o0,
			i1 => i19,
			o0 => Or259340_o0
		);
		Or259360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or259340_o0,
			i1 => i16,
			o0 => Or259360_o0
		);
		And259380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259360_o0,
			i1 => And2560_o0,
			o0 => And259380_o0
		);
		And259400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1280_o0,
			i1 => i5,
			o0 => And259400_o0
		);
		And259420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259400_o0,
			i1 => And211200_o0,
			o0 => And259420_o0
		);
		Or259440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259420_o0,
			i1 => And259380_o0,
			o0 => Or259440_o0
		);
		And259460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259440_o0,
			i1 => Not620_o0,
			o0 => And259460_o0
		);
		Or259480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259460_o0,
			i1 => And255900_o0,
			o0 => Or259480_o0
		);
		And259500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259480_o0,
			i1 => Nor29260_o0,
			o0 => And259500_o0
		);
		And259520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i13,
			i1 => Not540_o0,
			o0 => And259520_o0
		);
		And259540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259520_o0,
			i1 => And24040_o0,
			o0 => And259540_o0
		);
		Or259560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259540_o0,
			i1 => And259500_o0,
			o0 => Or259560_o0
		);
		And259580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259560_o0,
			i1 => i18,
			o0 => And259580_o0
		);
		Or259600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219920_o0,
			i1 => And219600_o0,
			o0 => Or259600_o0
		);
		And259620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259600_o0,
			i1 => Xor2960_o0,
			o0 => And259620_o0
		);
		And259640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28060_o0,
			i1 => i13,
			o0 => And259640_o0
		);
		Or259660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259640_o0,
			i1 => Nor29260_o0,
			o0 => Or259660_o0
		);
		And259680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259660_o0,
			i1 => Not7440_o0,
			o0 => And259680_o0
		);
		And259700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222020_o0,
			i1 => And219600_o0,
			o0 => And259700_o0
		);
		Or259720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259700_o0,
			i1 => And259680_o0,
			o0 => Or259720_o0
		);
		Or259740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or259720_o0,
			i1 => And259620_o0,
			o0 => Or259740_o0
		);
		And259760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259740_o0,
			i1 => And236120_o0,
			o0 => And259760_o0
		);
		Or259780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259760_o0,
			i1 => And259580_o0,
			o0 => Or259780_o0
		);
		And259800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259780_o0,
			i1 => i17,
			o0 => And259800_o0
		);
		And259820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => And25420_o0,
			o0 => And259820_o0
		);
		Or259840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And219920_o0,
			i1 => And219780_o0,
			o0 => Or259840_o0
		);
		Or259860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or259840_o0,
			i1 => And259820_o0,
			o0 => Or259860_o0
		);
		And259880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259860_o0,
			i1 => Not1500_o0,
			o0 => And259880_o0
		);
		And259900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2240_o0,
			i1 => i15,
			o0 => And259900_o0
		);
		And259920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259900_o0,
			i1 => Nor29260_o0,
			o0 => And259920_o0
		);
		Or259940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259920_o0,
			i1 => And259880_o0,
			o0 => Or259940_o0
		);
		And259960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or259940_o0,
			i1 => i16,
			o0 => And259960_o0
		);
		And259980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => Not620_o0,
			o0 => And259980_o0
		);
		Or260000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259980_o0,
			i1 => And228040_o0,
			o0 => Or260000_o0
		);
		And260020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260000_o0,
			i1 => And219600_o0,
			o0 => And260020_o0
		);
		And260040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => Not1280_o0,
			o0 => And260040_o0
		);
		Or260060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260040_o0,
			i1 => And222320_o0,
			o0 => Or260060_o0
		);
		Or260080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234780_o0,
			i1 => And219600_o0,
			o0 => Or260080_o0
		);
		And260100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260080_o0,
			i1 => Or260060_o0,
			o0 => And260100_o0
		);
		And260120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And237200_o0,
			i1 => Nor29260_o0,
			o0 => And260120_o0
		);
		And260140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259640_o0,
			i1 => And246660_o0,
			o0 => And260140_o0
		);
		Or260160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260140_o0,
			i1 => And260120_o0,
			o0 => Or260160_o0
		);
		Or260180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or260160_o0,
			i1 => And260100_o0,
			o0 => Or260180_o0
		);
		Or260200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or260180_o0,
			i1 => And260020_o0,
			o0 => Or260200_o0
		);
		Or260220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or260200_o0,
			i1 => And259960_o0,
			o0 => Or260220_o0
		);
		And260240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260220_o0,
			i1 => Not1040_o0,
			o0 => And260240_o0
		);
		Or260260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260240_o0,
			i1 => And223260_o0,
			o0 => Or260260_o0
		);
		And260280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260260_o0,
			i1 => And2560_o0,
			o0 => And260280_o0
		);
		Or260300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260280_o0,
			i1 => And259800_o0,
			o0 => Or260300_o0
		);
		And260320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260300_o0,
			i1 => i12,
			o0 => And260320_o0
		);
		And260340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225460_o0,
			i1 => Nor21840_o0,
			o0 => And260340_o0
		);
		Or260360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260340_o0,
			i1 => Or219480_o0,
			o0 => Or260360_o0
		);
		And260380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223260_o0,
			i1 => i40,
			o0 => And260380_o0
		);
		And260400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260380_o0,
			i1 => Nor232220_o0,
			o0 => And260400_o0
		);
		And260420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260400_o0,
			i1 => Or260360_o0,
			o0 => And260420_o0
		);
		Or260440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260420_o0,
			i1 => And260320_o0,
			o0 => Or260440_o0
		);
		And260460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260440_o0,
			i1 => Not140_o0,
			o0 => And260460_o0
		);
		And260480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => i12,
			o0 => And260480_o0
		);
		And260500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260480_o0,
			i1 => And227520_o0,
			o0 => And260500_o0
		);
		And260520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260500_o0,
			i1 => And23060_o0,
			o0 => And260520_o0
		);
		Or260540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260520_o0,
			i1 => And260460_o0,
			o0 => Or260540_o0
		);
		And260560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260540_o0,
			i1 => Not60_o0,
			o0 => And260560_o0
		);
		Or260580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260560_o0,
			i1 => And258100_o0,
			o0 => Or260580_o0
		);
		And260600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260580_o0,
			i1 => And258160_o0,
			o0 => And260600_o0
		);
		And260620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216560_o0,
			i1 => And213900_o0,
			o0 => And260620_o0
		);
		Or260640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260620_o0,
			i1 => And227100_o0,
			o0 => Or260640_o0
		);
		And260660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260640_o0,
			i1 => And26520_o0,
			o0 => And260660_o0
		);
		Nor260680 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i19,
			i1 => i14,
			o0 => Nor260680_o0
		);
		And260700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor260680_o0,
			i1 => And257940_o0,
			o0 => And260700_o0
		);
		And260720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260700_o0,
			i1 => And29860_o0,
			o0 => And260720_o0
		);
		Or260740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260720_o0,
			i1 => And260660_o0,
			o0 => Or260740_o0
		);
		And260760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260740_o0,
			i1 => Not540_o0,
			o0 => And260760_o0
		);
		And260780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And240360_o0,
			i1 => And213900_o0,
			o0 => And260780_o0
		);
		And260800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260780_o0,
			i1 => And247980_o0,
			o0 => And260800_o0
		);
		Or260820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260800_o0,
			i1 => And260760_o0,
			o0 => Or260820_o0
		);
		And260840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260820_o0,
			i1 => Not120_o0,
			o0 => And260840_o0
		);
		And260860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213900_o0,
			i1 => Not1500_o0,
			o0 => And260860_o0
		);
		And260880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260860_o0,
			i1 => And219060_o0,
			o0 => And260880_o0
		);
		And260900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260880_o0,
			i1 => And259180_o0,
			o0 => And260900_o0
		);
		Or260920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260900_o0,
			i1 => And260840_o0,
			o0 => Or260920_o0
		);
		And260940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or260920_o0,
			i1 => Not620_o0,
			o0 => And260940_o0
		);
		And260960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21140_o0,
			i1 => Not540_o0,
			o0 => And260960_o0
		);
		And260980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260960_o0,
			i1 => And246340_o0,
			o0 => And260980_o0
		);
		Or261000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And260980_o0,
			i1 => And260940_o0,
			o0 => Or261000_o0
		);
		And261020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261000_o0,
			i1 => Not1280_o0,
			o0 => And261020_o0
		);
		And261040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260960_o0,
			i1 => And246440_o0,
			o0 => And261040_o0
		);
		Or261060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261040_o0,
			i1 => And261020_o0,
			o0 => Or261060_o0
		);
		And261080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261060_o0,
			i1 => i18,
			o0 => And261080_o0
		);
		And261100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260960_o0,
			i1 => And257160_o0,
			o0 => And261100_o0
		);
		Or261120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261100_o0,
			i1 => And261080_o0,
			o0 => Or261120_o0
		);
		And261140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261120_o0,
			i1 => i17,
			o0 => And261140_o0
		);
		And261160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => Not180_o0,
			o0 => And261160_o0
		);
		And261180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261160_o0,
			i1 => And246660_o0,
			o0 => And261180_o0
		);
		Or261200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261180_o0,
			i1 => Or227080_o0,
			o0 => Or261200_o0
		);
		And261220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor236400_o0,
			i1 => i40,
			o0 => And261220_o0
		);
		And261240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261220_o0,
			i1 => Nor21140_o0,
			o0 => And261240_o0
		);
		And261260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261240_o0,
			i1 => Or261200_o0,
			o0 => And261260_o0
		);
		Or261280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261260_o0,
			i1 => And261140_o0,
			o0 => Or261280_o0
		);
		And261300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261280_o0,
			i1 => Not2080_o0,
			o0 => And261300_o0
		);
		And261320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor243420_o0,
			i1 => Not620_o0,
			o0 => And261320_o0
		);
		Or261340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or239480_o0,
			i1 => And217360_o0,
			o0 => Or261340_o0
		);
		Or261360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or261340_o0,
			i1 => And261320_o0,
			o0 => Or261360_o0
		);
		And261380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222800_o0,
			i1 => Nor21140_o0,
			o0 => And261380_o0
		);
		And261400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261380_o0,
			i1 => And257320_o0,
			o0 => And261400_o0
		);
		And261420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261400_o0,
			i1 => Or261360_o0,
			o0 => And261420_o0
		);
		Or261440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261420_o0,
			i1 => And261300_o0,
			o0 => Or261440_o0
		);
		And261460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261440_o0,
			i1 => Not160_o0,
			o0 => And261460_o0
		);
		And261480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210560_o0,
			i1 => i5,
			o0 => And261480_o0
		);
		And261500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217780_o0,
			i1 => Not540_o0,
			o0 => And261500_o0
		);
		Or261520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261500_o0,
			i1 => And261480_o0,
			o0 => Or261520_o0
		);
		And261540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261520_o0,
			i1 => Not7120_o0,
			o0 => And261540_o0
		);
		And261560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210740_o0,
			i1 => Not540_o0,
			o0 => And261560_o0
		);
		Or261580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261560_o0,
			i1 => And261540_o0,
			o0 => Or261580_o0
		);
		And261600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230240_o0,
			i1 => And23080_o0,
			o0 => And261600_o0
		);
		And261620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261600_o0,
			i1 => And26040_o0,
			o0 => And261620_o0
		);
		And261640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i27,
			i1 => i21,
			o0 => And261640_o0
		);
		And261660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261640_o0,
			i1 => Nor229280_o0,
			o0 => And261660_o0
		);
		And261680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261660_o0,
			i1 => And229320_o0,
			o0 => And261680_o0
		);
		And261700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261680_o0,
			i1 => And261620_o0,
			o0 => And261700_o0
		);
		And261720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261700_o0,
			i1 => Or261580_o0,
			o0 => And261720_o0
		);
		Or261740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261720_o0,
			i1 => And261460_o0,
			o0 => Or261740_o0
		);
		And261760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261740_o0,
			i1 => And256680_o0,
			o0 => And261760_o0
		);
		Or261780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And234180_o0,
			i1 => And218920_o0,
			o0 => Or261780_o0
		);
		And261800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261780_o0,
			i1 => i2,
			o0 => And261800_o0
		);
		And261820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or258220_o0,
			i1 => And29560_o0,
			o0 => And261820_o0
		);
		Or261840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261820_o0,
			i1 => And210540_o0,
			o0 => Or261840_o0
		);
		And261860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor235820_o0,
			i1 => i40,
			o0 => And261860_o0
		);
		And261880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261860_o0,
			i1 => Or261840_o0,
			o0 => And261880_o0
		);
		Or261900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261880_o0,
			i1 => And261800_o0,
			o0 => Or261900_o0
		);
		And261920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261900_o0,
			i1 => i27,
			o0 => And261920_o0
		);
		And261940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i21,
			o0 => And261940_o0
		);
		And261960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor235820_o0,
			i1 => i20,
			o0 => And261960_o0
		);
		And261980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261960_o0,
			i1 => And261940_o0,
			o0 => And261980_o0
		);
		Or262000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And261980_o0,
			i1 => And261920_o0,
			o0 => Or262000_o0
		);
		And262020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262000_o0,
			i1 => And26580_o0,
			o0 => And262020_o0
		);
		And262040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nand210020_o0,
			i1 => And24620_o0,
			o0 => And262040_o0
		);
		And262060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262040_o0,
			i1 => And261860_o0,
			o0 => And262060_o0
		);
		Or262080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262060_o0,
			i1 => And262020_o0,
			o0 => Or262080_o0
		);
		And262100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262080_o0,
			i1 => And213900_o0,
			o0 => And262100_o0
		);
		And262120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246180_o0,
			i1 => Nor235820_o0,
			o0 => And262120_o0
		);
		Or262140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262120_o0,
			i1 => And262100_o0,
			o0 => Or262140_o0
		);
		And262160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262140_o0,
			i1 => Not620_o0,
			o0 => And262160_o0
		);
		And262180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219620_o0,
			i1 => i12,
			o0 => And262180_o0
		);
		Or262200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262180_o0,
			i1 => And227100_o0,
			o0 => Or262200_o0
		);
		And262220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246320_o0,
			i1 => Nor235820_o0,
			o0 => And262220_o0
		);
		And262240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262220_o0,
			i1 => Or262200_o0,
			o0 => And262240_o0
		);
		Or262260 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262240_o0,
			i1 => And262160_o0,
			o0 => Or262260_o0
		);
		And262280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262260_o0,
			i1 => Not1500_o0,
			o0 => And262280_o0
		);
		And262300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213900_o0,
			i1 => And26600_o0,
			o0 => And262300_o0
		);
		Or262320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262300_o0,
			i1 => Or246500_o0,
			o0 => Or262320_o0
		);
		And262340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor235820_o0,
			i1 => And224580_o0,
			o0 => And262340_o0
		);
		And262360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262340_o0,
			i1 => Or262320_o0,
			o0 => And262360_o0
		);
		Or262380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262360_o0,
			i1 => And262280_o0,
			o0 => Or262380_o0
		);
		And262400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262380_o0,
			i1 => i17,
			o0 => And262400_o0
		);
		And262420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And251940_o0,
			i1 => And227100_o0,
			o0 => And262420_o0
		);
		Nor262440 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i37,
			i1 => i19,
			o0 => Nor262440_o0
		);
		And262460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor262440_o0,
			i1 => And25420_o0,
			o0 => And262460_o0
		);
		And262480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213900_o0,
			i1 => Nor212260_o0,
			o0 => And262480_o0
		);
		And262500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262480_o0,
			i1 => And262460_o0,
			o0 => And262500_o0
		);
		Or262520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262500_o0,
			i1 => And262420_o0,
			o0 => Or262520_o0
		);
		And262540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262520_o0,
			i1 => Not1280_o0,
			o0 => And262540_o0
		);
		Or262560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262540_o0,
			i1 => Or227080_o0,
			o0 => Or262560_o0
		);
		And262580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262560_o0,
			i1 => And235900_o0,
			o0 => And262580_o0
		);
		Or262600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262580_o0,
			i1 => And262400_o0,
			o0 => Or262600_o0
		);
		And262620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262600_o0,
			i1 => Not2080_o0,
			o0 => And262620_o0
		);
		Or262640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And227280_o0,
			i1 => And210440_o0,
			o0 => Or262640_o0
		);
		Or262660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or262640_o0,
			i1 => And228200_o0,
			o0 => Or262660_o0
		);
		And262680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262660_o0,
			i1 => And22560_o0,
			o0 => And262680_o0
		);
		And262700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24000_o0,
			i1 => And21300_o0,
			o0 => And262700_o0
		);
		And262720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262700_o0,
			i1 => And212880_o0,
			o0 => And262720_o0
		);
		And262740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262720_o0,
			i1 => And212280_o0,
			o0 => And262740_o0
		);
		And262760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246960_o0,
			i1 => And21120_o0,
			o0 => And262760_o0
		);
		Or262780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262760_o0,
			i1 => And262740_o0,
			o0 => Or262780_o0
		);
		Or262800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or262780_o0,
			i1 => And262680_o0,
			o0 => Or262800_o0
		);
		And262820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i13,
			o0 => And262820_o0
		);
		And262840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262820_o0,
			i1 => Nor235820_o0,
			o0 => And262840_o0
		);
		And262860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And262840_o0,
			i1 => Or262800_o0,
			o0 => And262860_o0
		);
		Or262880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262860_o0,
			i1 => And262620_o0,
			o0 => Or262880_o0
		);
		And262900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262880_o0,
			i1 => Not160_o0,
			o0 => And262900_o0
		);
		And262920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And214880_o0,
			i1 => Not120_o0,
			o0 => And262920_o0
		);
		Or262940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And262920_o0,
			i1 => And262900_o0,
			o0 => Or262940_o0
		);
		And262960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or262940_o0,
			i1 => Not140_o0,
			o0 => And262960_o0
		);
		And262980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And230000_o0,
			i1 => i4,
			o0 => And262980_o0
		);
		And263000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215860_o0,
			i1 => i22,
			o0 => And263000_o0
		);
		And263020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254820_o0,
			i1 => i26,
			o0 => And263020_o0
		);
		And263040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263020_o0,
			i1 => And263000_o0,
			o0 => And263040_o0
		);
		Or263060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263040_o0,
			i1 => And262980_o0,
			o0 => Or263060_o0
		);
		And263080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263060_o0,
			i1 => i27,
			o0 => And263080_o0
		);
		And263100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254820_o0,
			i1 => And256740_o0,
			o0 => And263100_o0
		);
		And263120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263100_o0,
			i1 => And263000_o0,
			o0 => And263120_o0
		);
		Or263140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263120_o0,
			i1 => And263080_o0,
			o0 => Or263140_o0
		);
		And263160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26040_o0,
			i1 => And23080_o0,
			o0 => And263160_o0
		);
		And263180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263160_o0,
			i1 => And218980_o0,
			o0 => And263180_o0
		);
		And263200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263180_o0,
			i1 => And248260_o0,
			o0 => And263200_o0
		);
		And263220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263200_o0,
			i1 => Or263140_o0,
			o0 => And263220_o0
		);
		Or263240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263220_o0,
			i1 => And262960_o0,
			o0 => Or263240_o0
		);
		Nor263260 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i9,
			o0 => Nor263260_o0
		);
		And263280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor263260_o0,
			i1 => Nor23600_o0,
			o0 => And263280_o0
		);
		And263300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263280_o0,
			i1 => Or263240_o0,
			o0 => And263300_o0
		);
		Or263320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263300_o0,
			i1 => i9,
			o0 => Or263320_o0
		);
		And263340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263320_o0,
			i1 => Not24960_o0,
			o0 => And263340_o0
		);
		And263360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			i1 => i9,
			o0 => And263360_o0
		);
		Or263380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263360_o0,
			i1 => And263340_o0,
			o0 => Or263380_o0
		);
		And263400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263380_o0,
			i1 => Not12120_o0,
			o0 => And263400_o0
		);
		Or263420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263400_o0,
			i1 => And220460_o0,
			o0 => Or263420_o0
		);
		And263440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263420_o0,
			i1 => Not12100_o0,
			o0 => And263440_o0
		);
		And263460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => Not1280_o0,
			o0 => And263460_o0
		);
		And263480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215060_o0,
			i1 => i16,
			o0 => And263480_o0
		);
		Or263500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263480_o0,
			i1 => And263460_o0,
			o0 => Or263500_o0
		);
		And263520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263500_o0,
			i1 => Not620_o0,
			o0 => And263520_o0
		);
		Or263540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263520_o0,
			i1 => And246800_o0,
			o0 => Or263540_o0
		);
		And263560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263540_o0,
			i1 => Not1040_o0,
			o0 => And263560_o0
		);
		And263580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => i16,
			o0 => And263580_o0
		);
		And263600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263580_o0,
			i1 => Not620_o0,
			o0 => And263600_o0
		);
		Or263620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263600_o0,
			i1 => And263560_o0,
			o0 => Or263620_o0
		);
		And263640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263620_o0,
			i1 => i13,
			o0 => And263640_o0
		);
		And263660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => i16,
			o0 => And263660_o0
		);
		Or263680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263660_o0,
			i1 => And254980_o0,
			o0 => Or263680_o0
		);
		Or263700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or263680_o0,
			i1 => Not2080_o0,
			o0 => Or263700_o0
		);
		Or263720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or263700_o0,
			i1 => And263640_o0,
			o0 => Or263720_o0
		);
		And263740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263720_o0,
			i1 => i14,
			o0 => And263740_o0
		);
		Or263760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217340_o0,
			i1 => And22380_o0,
			o0 => Or263760_o0
		);
		And263780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263760_o0,
			i1 => i15,
			o0 => And263780_o0
		);
		And263800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22300_o0,
			i1 => Not1080_o0,
			o0 => And263800_o0
		);
		And263820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263800_o0,
			i1 => Or217020_o0,
			o0 => And263820_o0
		);
		Or263840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263820_o0,
			i1 => And263780_o0,
			o0 => Or263840_o0
		);
		And263860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263840_o0,
			i1 => i16,
			o0 => And263860_o0
		);
		And263880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228740_o0,
			i1 => And21300_o0,
			o0 => And263880_o0
		);
		Or263900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263880_o0,
			i1 => And263860_o0,
			o0 => Or263900_o0
		);
		And263920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263900_o0,
			i1 => Nor29260_o0,
			o0 => And263920_o0
		);
		Or263940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263920_o0,
			i1 => And263740_o0,
			o0 => Or263940_o0
		);
		And263960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or263940_o0,
			i1 => i12,
			o0 => And263960_o0
		);
		And263980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => Nor2220_o0,
			o0 => And263980_o0
		);
		And264000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213700_o0,
			i1 => i13,
			o0 => And264000_o0
		);
		And264020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => Not1080_o0,
			o0 => And264020_o0
		);
		Or264040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264020_o0,
			i1 => And264000_o0,
			o0 => Or264040_o0
		);
		Or264060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264040_o0,
			i1 => And263980_o0,
			o0 => Or264060_o0
		);
		And264080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264060_o0,
			i1 => i12,
			o0 => And264080_o0
		);
		And264100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => i14,
			o0 => And264100_o0
		);
		And264120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And264100_o0,
			i1 => Nor224000_o0,
			o0 => And264120_o0
		);
		Or264140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264120_o0,
			i1 => And264080_o0,
			o0 => Or264140_o0
		);
		And264160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264140_o0,
			i1 => i15,
			o0 => And264160_o0
		);
		And264180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or235220_o0,
			i1 => i12,
			o0 => And264180_o0
		);
		And264200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223260_o0,
			i1 => Not180_o0,
			o0 => And264200_o0
		);
		Or264220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264200_o0,
			i1 => And264180_o0,
			o0 => Or264220_o0
		);
		And264240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264220_o0,
			i1 => i17,
			o0 => And264240_o0
		);
		And264260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => i14,
			o0 => And264260_o0
		);
		And264280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And264260_o0,
			i1 => Nor224000_o0,
			o0 => And264280_o0
		);
		Or264300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264280_o0,
			i1 => And264240_o0,
			o0 => Or264300_o0
		);
		Or264320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264300_o0,
			i1 => And264160_o0,
			o0 => Or264320_o0
		);
		And264340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264320_o0,
			i1 => Xor2960_o0,
			o0 => And264340_o0
		);
		And264360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228580_o0,
			i1 => Nor29260_o0,
			o0 => And264360_o0
		);
		Nor264380 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i17,
			i1 => i15,
			o0 => Nor264380_o0
		);
		And264400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => Nor264380_o0,
			o0 => And264400_o0
		);
		Or264420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264400_o0,
			i1 => And264360_o0,
			o0 => Or264420_o0
		);
		And264440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264420_o0,
			i1 => i12,
			o0 => And264440_o0
		);
		Or264460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And259640_o0,
			i1 => And234780_o0,
			o0 => Or264460_o0
		);
		And264480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264460_o0,
			i1 => i12,
			o0 => And264480_o0
		);
		And264500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor224000_o0,
			i1 => And28060_o0,
			o0 => And264500_o0
		);
		And264520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22300_o0,
			i1 => i14,
			o0 => And264520_o0
		);
		And264540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And264520_o0,
			i1 => Nor224000_o0,
			o0 => And264540_o0
		);
		Or264560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264540_o0,
			i1 => And264500_o0,
			o0 => Or264560_o0
		);
		Or264580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264560_o0,
			i1 => And264480_o0,
			o0 => Or264580_o0
		);
		Or264600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264580_o0,
			i1 => And264440_o0,
			o0 => Or264600_o0
		);
		And264620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264600_o0,
			i1 => Or260060_o0,
			o0 => And264620_o0
		);
		And264640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not28160_o0,
			i1 => And21060_o0,
			o0 => And264640_o0
		);
		Or264660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264640_o0,
			i1 => And254980_o0,
			o0 => Or264660_o0
		);
		And264680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264660_o0,
			i1 => Not620_o0,
			o0 => And264680_o0
		);
		Or264700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And263660_o0,
			i1 => And254620_o0,
			o0 => Or264700_o0
		);
		And264720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264700_o0,
			i1 => i15,
			o0 => And264720_o0
		);
		And264740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21100_o0,
			i1 => And2640_o0,
			o0 => And264740_o0
		);
		Or264760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264740_o0,
			i1 => And264720_o0,
			o0 => Or264760_o0
		);
		Or264780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264760_o0,
			i1 => And264680_o0,
			o0 => Or264780_o0
		);
		And264800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor224000_o0,
			i1 => i14,
			o0 => And264800_o0
		);
		And264820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And264800_o0,
			i1 => Or264780_o0,
			o0 => And264820_o0
		);
		Or264840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264820_o0,
			i1 => And264620_o0,
			o0 => Or264840_o0
		);
		Or264860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264840_o0,
			i1 => And264340_o0,
			o0 => Or264860_o0
		);
		Or264880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or264860_o0,
			i1 => And263960_o0,
			o0 => Or264880_o0
		);
		And264900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264880_o0,
			i1 => And26520_o0,
			o0 => And264900_o0
		);
		Or264920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264900_o0,
			i1 => And257980_o0,
			o0 => Or264920_o0
		);
		And264940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or264920_o0,
			i1 => Not60_o0,
			o0 => And264940_o0
		);
		And264960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260480_o0,
			i1 => And26760_o0,
			o0 => And264960_o0
		);
		And264980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And264960_o0,
			i1 => And23060_o0,
			o0 => And264980_o0
		);
		Or265000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And264980_o0,
			i1 => And264940_o0,
			o0 => Or265000_o0
		);
		And265020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213260_o0,
			i1 => Nor22060_o0,
			o0 => And265020_o0
		);
		And265040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265020_o0,
			i1 => And23340_o0,
			o0 => And265040_o0
		);
		And265060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265040_o0,
			i1 => Or265000_o0,
			o0 => And265060_o0
		);
		And265080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or24600_o0,
			i1 => Xor2960_o0,
			o0 => And265080_o0
		);
		And265100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25280_o0,
			i1 => Not540_o0,
			o0 => And265100_o0
		);
		And265120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265100_o0,
			i1 => And25040_o0,
			o0 => And265120_o0
		);
		Or265140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265120_o0,
			i1 => And265080_o0,
			o0 => Or265140_o0
		);
		And265160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265140_o0,
			i1 => i1,
			o0 => And265160_o0
		);
		And265180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210400_o0,
			i1 => Not160_o0,
			o0 => And265180_o0
		);
		And265200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22060_o0,
			i1 => Not140_o0,
			o0 => And265200_o0
		);
		And265220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265200_o0,
			i1 => And265180_o0,
			o0 => And265220_o0
		);
		And265240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or25060_o0,
			i1 => Not100_o0,
			o0 => And265240_o0
		);
		And265260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224460_o0,
			i1 => Nor22600_o0,
			o0 => And265260_o0
		);
		And265280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i1,
			o0 => And265280_o0
		);
		And265300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not540_o0,
			o0 => And265300_o0
		);
		And265320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265300_o0,
			i1 => And265280_o0,
			o0 => And265320_o0
		);
		And265340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265320_o0,
			i1 => Nor21140_o0,
			o0 => And265340_o0
		);
		Or265360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265340_o0,
			i1 => And265260_o0,
			o0 => Or265360_o0
		);
		Or265380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or265360_o0,
			i1 => And265240_o0,
			o0 => Or265380_o0
		);
		Or265400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or265380_o0,
			i1 => And265220_o0,
			o0 => Or265400_o0
		);
		Or265420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or265400_o0,
			i1 => And265160_o0,
			o0 => Or265420_o0
		);
		And265440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265420_o0,
			i1 => And27500_o0,
			o0 => And265440_o0
		);
		And265460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25020_o0,
			i1 => Nor22060_o0,
			o0 => And265460_o0
		);
		Or265480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265460_o0,
			i1 => Or26100_o0,
			o0 => Or265480_o0
		);
		Or265500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or265480_o0,
			i1 => And265220_o0,
			o0 => Or265500_o0
		);
		And265520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26120_o0,
			i1 => And2640_o0,
			o0 => And265520_o0
		);
		And265540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265520_o0,
			i1 => Or265500_o0,
			o0 => And265540_o0
		);
		Or265560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265540_o0,
			i1 => And265440_o0,
			o0 => Or265560_o0
		);
		And265580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265560_o0,
			i1 => Not60_o0,
			o0 => And265580_o0
		);
		And265600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or224860_o0,
			i1 => And211740_o0,
			o0 => And265600_o0
		);
		Or265620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265600_o0,
			i1 => And265580_o0,
			o0 => Or265620_o0
		);
		And265640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23280_o0,
			i1 => And23020_o0,
			o0 => And265640_o0
		);
		And265660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265640_o0,
			i1 => And215720_o0,
			o0 => And265660_o0
		);
		And265680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265660_o0,
			i1 => Or265620_o0,
			o0 => And265680_o0
		);
		And265700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2980_o0,
			i1 => Not180_o0,
			o0 => And265700_o0
		);
		And265720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265700_o0,
			i1 => i4,
			o0 => And265720_o0
		);
		And265740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25840_o0,
			i1 => Not160_o0,
			o0 => And265740_o0
		);
		Or265760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265740_o0,
			i1 => And265720_o0,
			o0 => Or265760_o0
		);
		And265780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265760_o0,
			i1 => Not140_o0,
			o0 => And265780_o0
		);
		And265800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265700_o0,
			i1 => i3,
			o0 => And265800_o0
		);
		Or265820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265800_o0,
			i1 => And265780_o0,
			o0 => Or265820_o0
		);
		And265840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265820_o0,
			i1 => Not120_o0,
			o0 => And265840_o0
		);
		And265860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265700_o0,
			i1 => i2,
			o0 => And265860_o0
		);
		Or265880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265860_o0,
			i1 => And265840_o0,
			o0 => Or265880_o0
		);
		And265900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265880_o0,
			i1 => Not100_o0,
			o0 => And265900_o0
		);
		And265920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265700_o0,
			i1 => i1,
			o0 => And265920_o0
		);
		Or265940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And265920_o0,
			i1 => And265900_o0,
			o0 => Or265940_o0
		);
		And265960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or265940_o0,
			i1 => Not540_o0,
			o0 => And265960_o0
		);
		And265980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24280_o0,
			i1 => Nor2220_o0,
			o0 => And265980_o0
		);
		And266000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And265980_o0,
			i1 => Xor2960_o0,
			o0 => And266000_o0
		);
		And266020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266000_o0,
			i1 => Or265480_o0,
			o0 => And266020_o0
		);
		Or266040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266020_o0,
			i1 => And265960_o0,
			o0 => Or266040_o0
		);
		And266060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266040_o0,
			i1 => i15,
			o0 => And266060_o0
		);
		Or266080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i3,
			o0 => Or266080_o0
		);
		And266100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266080_o0,
			i1 => And21640_o0,
			o0 => And266100_o0
		);
		And266120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215440_o0,
			i1 => Nor22600_o0,
			o0 => And266120_o0
		);
		Or266140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266120_o0,
			i1 => And266100_o0,
			o0 => Or266140_o0
		);
		And266160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24880_o0,
			i1 => i19,
			o0 => And266160_o0
		);
		And266180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266160_o0,
			i1 => Or266140_o0,
			o0 => And266180_o0
		);
		And266200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25840_o0,
			i1 => Nor22600_o0,
			o0 => And266200_o0
		);
		Or266220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266200_o0,
			i1 => And266180_o0,
			o0 => Or266220_o0
		);
		And266240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266220_o0,
			i1 => Not120_o0,
			o0 => And266240_o0
		);
		And266260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25940_o0,
			i1 => Not180_o0,
			o0 => And266260_o0
		);
		And266280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266260_o0,
			i1 => i2,
			o0 => And266280_o0
		);
		Or266300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266280_o0,
			i1 => And266240_o0,
			o0 => Or266300_o0
		);
		And266320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266300_o0,
			i1 => Not100_o0,
			o0 => And266320_o0
		);
		And266340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266260_o0,
			i1 => i1,
			o0 => And266340_o0
		);
		Or266360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266340_o0,
			i1 => And266320_o0,
			o0 => Or266360_o0
		);
		And266380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266360_o0,
			i1 => Not540_o0,
			o0 => And266380_o0
		);
		And266400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And210420_o0,
			i1 => And2240_o0,
			o0 => And266400_o0
		);
		And266420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266400_o0,
			i1 => And24280_o0,
			o0 => And266420_o0
		);
		And266440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266420_o0,
			i1 => Or265480_o0,
			o0 => And266440_o0
		);
		Or266460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266440_o0,
			i1 => And266380_o0,
			o0 => Or266460_o0
		);
		And266480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266460_o0,
			i1 => Not620_o0,
			o0 => And266480_o0
		);
		Or266500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266480_o0,
			i1 => And266060_o0,
			o0 => Or266500_o0
		);
		And266520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266500_o0,
			i1 => Not60_o0,
			o0 => And266520_o0
		);
		Or266540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266520_o0,
			i1 => And29000_o0,
			o0 => Or266540_o0
		);
		And266560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266540_o0,
			i1 => i13,
			o0 => And266560_o0
		);
		Nor266580 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor228140_o0,
			i1 => i16,
			o0 => Nor266580_o0
		);
		Or266600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Nor266580_o0,
			i1 => And222320_o0,
			o0 => Or266600_o0
		);
		And266620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266600_o0,
			i1 => Not620_o0,
			o0 => And266620_o0
		);
		Or266640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266620_o0,
			i1 => And254560_o0,
			o0 => Or266640_o0
		);
		And266660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266640_o0,
			i1 => i17,
			o0 => And266660_o0
		);
		And266680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And218580_o0,
			i1 => And21300_o0,
			o0 => And266680_o0
		);
		Or266700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266680_o0,
			i1 => And266660_o0,
			o0 => Or266700_o0
		);
		And266720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266700_o0,
			i1 => And2560_o0,
			o0 => And266720_o0
		);
		Or266740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266720_o0,
			i1 => And21880_o0,
			o0 => Or266740_o0
		);
		And266760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266740_o0,
			i1 => Not140_o0,
			o0 => And266760_o0
		);
		Or266780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266760_o0,
			i1 => And22020_o0,
			o0 => Or266780_o0
		);
		And266800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266780_o0,
			i1 => Not60_o0,
			o0 => And266800_o0
		);
		And266820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And26760_o0,
			i1 => Nor21980_o0,
			o0 => And266820_o0
		);
		And266840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266820_o0,
			i1 => And21960_o0,
			o0 => And266840_o0
		);
		Or266860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266840_o0,
			i1 => And266800_o0,
			o0 => Or266860_o0
		);
		And266880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266860_o0,
			i1 => And22140_o0,
			o0 => And266880_o0
		);
		Or266900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And266880_o0,
			i1 => And266560_o0,
			o0 => Or266900_o0
		);
		And266920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or266900_o0,
			i1 => Not80_o0,
			o0 => And266920_o0
		);
		Or266940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And217360_o0,
			i1 => And22800_o0,
			o0 => Or266940_o0
		);
		Or266960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or266940_o0,
			i1 => Not2080_o0,
			o0 => Or266960_o0
		);
		And266980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22560_o0,
			i1 => Nor21140_o0,
			o0 => And266980_o0
		);
		And267000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And266980_o0,
			i1 => Nor23600_o0,
			o0 => And267000_o0
		);
		And267020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267000_o0,
			i1 => And216700_o0,
			o0 => And267020_o0
		);
		And267040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267020_o0,
			i1 => Or266960_o0,
			o0 => And267040_o0
		);
		Or267060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267040_o0,
			i1 => And266920_o0,
			o0 => Or267060_o0
		);
		And267080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267060_o0,
			i1 => And23360_o0,
			o0 => And267080_o0
		);
		And267100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or215920_o0,
			i1 => i1,
			o0 => And267100_o0
		);
		And267120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor25100_o0,
			i1 => Xor2960_o0,
			o0 => And267120_o0
		);
		And267140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267120_o0,
			i1 => Or210400_o0,
			o0 => And267140_o0
		);
		Or267160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267140_o0,
			i1 => And267100_o0,
			o0 => Or267160_o0
		);
		And267180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267160_o0,
			i1 => Nor24000_o0,
			o0 => And267180_o0
		);
		And267200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor25100_o0,
			i1 => Not540_o0,
			o0 => And267200_o0
		);
		And267220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267200_o0,
			i1 => And24060_o0,
			o0 => And267220_o0
		);
		Or267240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267220_o0,
			i1 => And267180_o0,
			o0 => Or267240_o0
		);
		And267260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267240_o0,
			i1 => i15,
			o0 => And267260_o0
		);
		Or267280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Not80_o0,
			i1 => i12,
			o0 => Or267280_o0
		);
		And267300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267280_o0,
			i1 => Not1500_o0,
			o0 => And267300_o0
		);
		And267320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246260_o0,
			i1 => Not180_o0,
			o0 => And267320_o0
		);
		Or267340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267320_o0,
			i1 => And267300_o0,
			o0 => Or267340_o0
		);
		And267360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267340_o0,
			i1 => i16,
			o0 => And267360_o0
		);
		And267380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215880_o0,
			i1 => And22560_o0,
			o0 => And267380_o0
		);
		Or267400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267380_o0,
			i1 => And267360_o0,
			o0 => Or267400_o0
		);
		And267420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21980_o0,
			i1 => i40,
			o0 => And267420_o0
		);
		And267440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267420_o0,
			i1 => Nor25100_o0,
			o0 => And267440_o0
		);
		And267460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267440_o0,
			i1 => Or267400_o0,
			o0 => And267460_o0
		);
		Or267480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267460_o0,
			i1 => And267260_o0,
			o0 => Or267480_o0
		);
		And267500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267480_o0,
			i1 => Not1080_o0,
			o0 => And267500_o0
		);
		And267520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222800_o0,
			i1 => And28060_o0,
			o0 => And267520_o0
		);
		And267540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor25100_o0,
			i1 => And24180_o0,
			o0 => And267540_o0
		);
		And267560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267540_o0,
			i1 => And267520_o0,
			o0 => And267560_o0
		);
		Or267580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267560_o0,
			i1 => And267500_o0,
			o0 => Or267580_o0
		);
		And267600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267580_o0,
			i1 => Not1040_o0,
			o0 => And267600_o0
		);
		Nor267620 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i12,
			o0 => Nor267620_o0
		);
		And267640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor267620_o0,
			i1 => And2260_o0,
			o0 => And267640_o0
		);
		Or267660 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267640_o0,
			i1 => i12,
			o0 => Or267660_o0
		);
		And267680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267660_o0,
			i1 => i15,
			o0 => And267680_o0
		);
		And267700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => Not180_o0,
			o0 => And267700_o0
		);
		And267720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267700_o0,
			i1 => And2260_o0,
			o0 => And267720_o0
		);
		Or267740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267720_o0,
			i1 => And267680_o0,
			o0 => Or267740_o0
		);
		And267760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267740_o0,
			i1 => Not80_o0,
			o0 => And267760_o0
		);
		And267780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22560_o0,
			i1 => Nor21840_o0,
			o0 => And267780_o0
		);
		And267800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267780_o0,
			i1 => And214100_o0,
			o0 => And267800_o0
		);
		Or267820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267800_o0,
			i1 => And267760_o0,
			o0 => Or267820_o0
		);
		And267840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267820_o0,
			i1 => And2560_o0,
			o0 => And267840_o0
		);
		And267860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => And24280_o0,
			o0 => And267860_o0
		);
		And267880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And267860_o0,
			i1 => And266400_o0,
			o0 => And267880_o0
		);
		Or267900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267880_o0,
			i1 => And267840_o0,
			o0 => Or267900_o0
		);
		And267920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267900_o0,
			i1 => Nor25100_o0,
			o0 => And267920_o0
		);
		Or267940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And267920_o0,
			i1 => And267600_o0,
			o0 => Or267940_o0
		);
		And267960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267940_o0,
			i1 => i13,
			o0 => And267960_o0
		);
		Or267980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21240_o0,
			i1 => And2260_o0,
			o0 => Or267980_o0
		);
		And268000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or267980_o0,
			i1 => Not620_o0,
			o0 => And268000_o0
		);
		And268020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or244200_o0,
			i1 => i15,
			o0 => And268020_o0
		);
		Or268040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268020_o0,
			i1 => And268000_o0,
			o0 => Or268040_o0
		);
		And268060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268040_o0,
			i1 => Not1280_o0,
			o0 => And268060_o0
		);
		Or268080 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268060_o0,
			i1 => And21760_o0,
			o0 => Or268080_o0
		);
		And268100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268080_o0,
			i1 => Not80_o0,
			o0 => And268100_o0
		);
		And268120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor252020_o0,
			i1 => And21820_o0,
			o0 => And268120_o0
		);
		Or268140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268120_o0,
			i1 => i14,
			o0 => Or268140_o0
		);
		Or268160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or268140_o0,
			i1 => And268100_o0,
			o0 => Or268160_o0
		);
		And268180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268160_o0,
			i1 => And2560_o0,
			o0 => And268180_o0
		);
		And268200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => i5,
			o0 => And268200_o0
		);
		And268220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268200_o0,
			i1 => And21960_o0,
			o0 => And268220_o0
		);
		Or268240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268220_o0,
			i1 => And268180_o0,
			o0 => Or268240_o0
		);
		And268260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor25100_o0,
			i1 => And23080_o0,
			o0 => And268260_o0
		);
		And268280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268260_o0,
			i1 => Or268240_o0,
			o0 => And268280_o0
		);
		Or268300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268280_o0,
			i1 => And267960_o0,
			o0 => Or268300_o0
		);
		And268320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268300_o0,
			i1 => Not60_o0,
			o0 => And268320_o0
		);
		And268340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239120_o0,
			i1 => i4,
			o0 => And268340_o0
		);
		Or268360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268340_o0,
			i1 => And211700_o0,
			o0 => Or268360_o0
		);
		And268380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23180_o0,
			i1 => Not80_o0,
			o0 => And268380_o0
		);
		And268400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268380_o0,
			i1 => Or268360_o0,
			o0 => And268400_o0
		);
		Or268420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268400_o0,
			i1 => And268320_o0,
			o0 => Or268420_o0
		);
		And268440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268420_o0,
			i1 => Not140_o0,
			o0 => And268440_o0
		);
		And268460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And239120_o0,
			i1 => i0,
			o0 => And268460_o0
		);
		And268480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And254700_o0,
			i1 => Nor211040_o0,
			o0 => And268480_o0
		);
		And268500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268480_o0,
			i1 => And21960_o0,
			o0 => And268500_o0
		);
		Or268520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268500_o0,
			i1 => And268460_o0,
			o0 => Or268520_o0
		);
		And268540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227520_o0,
			i1 => Not80_o0,
			o0 => And268540_o0
		);
		And268560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268540_o0,
			i1 => Nor25100_o0,
			o0 => And268560_o0
		);
		And268580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268560_o0,
			i1 => Or268520_o0,
			o0 => And268580_o0
		);
		Or268600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268580_o0,
			i1 => And268440_o0,
			o0 => Or268600_o0
		);
		And268620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214980_o0,
			i1 => Nor212700_o0,
			o0 => And268620_o0
		);
		And268640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268620_o0,
			i1 => Nor248660_o0,
			o0 => And268640_o0
		);
		And268660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268640_o0,
			i1 => Or268600_o0,
			o0 => And268660_o0
		);
		And268680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or28520_o0,
			i1 => And23020_o0,
			o0 => And268680_o0
		);
		And268700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25600_o0,
			i1 => Not620_o0,
			o0 => And268700_o0
		);
		And268720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268700_o0,
			i1 => And23100_o0,
			o0 => And268720_o0
		);
		Or268740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268720_o0,
			i1 => And268680_o0,
			o0 => Or268740_o0
		);
		And268760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268740_o0,
			i1 => Not1040_o0,
			o0 => And268760_o0
		);
		And268780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223240_o0,
			i1 => And21300_o0,
			o0 => And268780_o0
		);
		And268800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268780_o0,
			i1 => And23100_o0,
			o0 => And268800_o0
		);
		Or268820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268800_o0,
			i1 => And268760_o0,
			o0 => Or268820_o0
		);
		And268840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268820_o0,
			i1 => Not1500_o0,
			o0 => And268840_o0
		);
		And268860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24280_o0,
			i1 => i13,
			o0 => And268860_o0
		);
		And268880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268860_o0,
			i1 => And231440_o0,
			o0 => And268880_o0
		);
		Or268900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268880_o0,
			i1 => And268840_o0,
			o0 => Or268900_o0
		);
		And268920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or268900_o0,
			i1 => Not160_o0,
			o0 => And268920_o0
		);
		And268940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And22800_o0,
			o0 => And268940_o0
		);
		And268960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268940_o0,
			i1 => Not7440_o0,
			o0 => And268960_o0
		);
		And268980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268960_o0,
			i1 => i4,
			o0 => And268980_o0
		);
		Or269000 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And268980_o0,
			i1 => And268920_o0,
			o0 => Or269000_o0
		);
		And269020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269000_o0,
			i1 => Not140_o0,
			o0 => And269020_o0
		);
		And269040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268960_o0,
			i1 => i3,
			o0 => And269040_o0
		);
		Or269060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269040_o0,
			i1 => And269020_o0,
			o0 => Or269060_o0
		);
		And269080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269060_o0,
			i1 => Not120_o0,
			o0 => And269080_o0
		);
		And269100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And268960_o0,
			i1 => i2,
			o0 => And269100_o0
		);
		Or269120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269100_o0,
			i1 => And269080_o0,
			o0 => Or269120_o0
		);
		And269140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269120_o0,
			i1 => Not1080_o0,
			o0 => And269140_o0
		);
		And269160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And25600_o0,
			i1 => And22940_o0,
			o0 => And269160_o0
		);
		Or269180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269160_o0,
			i1 => And216280_o0,
			o0 => Or269180_o0
		);
		And269200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225680_o0,
			i1 => And214100_o0,
			o0 => And269200_o0
		);
		Nor269220 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i12,
			i1 => i4,
			o0 => Nor269220_o0
		);
		And269240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor269220_o0,
			i1 => Nor21140_o0,
			o0 => And269240_o0
		);
		And269260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269240_o0,
			i1 => And269200_o0,
			o0 => And269260_o0
		);
		And269280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269260_o0,
			i1 => Or269180_o0,
			o0 => And269280_o0
		);
		Or269300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269280_o0,
			i1 => And269140_o0,
			o0 => Or269300_o0
		);
		And269320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269300_o0,
			i1 => Not60_o0,
			o0 => And269320_o0
		);
		Xor269340 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i3,
			o0 => Xor269340_o0
		);
		And269360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor269220_o0,
			i1 => And22480_o0,
			o0 => And269360_o0
		);
		And269380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269360_o0,
			i1 => And237440_o0,
			o0 => And269380_o0
		);
		And269400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269380_o0,
			i1 => Xor269340_o0,
			o0 => And269400_o0
		);
		And269420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269400_o0,
			i1 => Or22840_o0,
			o0 => And269420_o0
		);
		Or269440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269420_o0,
			i1 => And269320_o0,
			o0 => Or269440_o0
		);
		And269460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269440_o0,
			i1 => Not100_o0,
			o0 => And269460_o0
		);
		Nor269480 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor25220_o0,
			i1 => i5,
			o0 => Nor269480_o0
		);
		And269500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215820_o0,
			i1 => i5,
			o0 => And269500_o0
		);
		Or269520 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269500_o0,
			i1 => Nor269480_o0,
			o0 => Or269520_o0
		);
		And269540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225320_o0,
			i1 => Nor2220_o0,
			o0 => And269540_o0
		);
		And269560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor269220_o0,
			i1 => And224460_o0,
			o0 => And269560_o0
		);
		And269580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269560_o0,
			i1 => Nor237580_o0,
			o0 => And269580_o0
		);
		And269600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269580_o0,
			i1 => And269540_o0,
			o0 => And269600_o0
		);
		And269620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269600_o0,
			i1 => Or269520_o0,
			o0 => And269620_o0
		);
		Or269640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269620_o0,
			i1 => And269460_o0,
			o0 => Or269640_o0
		);
		And269660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269640_o0,
			i1 => Not80_o0,
			o0 => And269660_o0
		);
		And269680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222800_o0,
			i1 => And219600_o0,
			o0 => And269680_o0
		);
		And269700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269680_o0,
			i1 => And22620_o0,
			o0 => And269700_o0
		);
		And269720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And222120_o0,
			i1 => Nor2220_o0,
			o0 => And269720_o0
		);
		And269740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => Not60_o0,
			o0 => And269740_o0
		);
		And269760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269740_o0,
			i1 => And269720_o0,
			o0 => And269760_o0
		);
		And269780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269760_o0,
			i1 => And269700_o0,
			o0 => And269780_o0
		);
		Or269800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269780_o0,
			i1 => And269660_o0,
			o0 => Or269800_o0
		);
		And269820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269800_o0,
			i1 => And23360_o0,
			o0 => And269820_o0
		);
		And269840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And217280_o0,
			i1 => And23080_o0,
			o0 => And269840_o0
		);
		And269860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21060_o0,
			i1 => i15,
			o0 => And269860_o0
		);
		And269880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269860_o0,
			i1 => And23020_o0,
			o0 => And269880_o0
		);
		Or269900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269880_o0,
			i1 => And269840_o0,
			o0 => Or269900_o0
		);
		And269920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or269900_o0,
			i1 => i5,
			o0 => And269920_o0
		);
		And269940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => And21940_o0,
			o0 => And269940_o0
		);
		And269960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And21060_o0,
			o0 => And269960_o0
		);
		Or269980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And269960_o0,
			i1 => And269940_o0,
			o0 => Or269980_o0
		);
		And270000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22940_o0,
			i1 => i40,
			o0 => And270000_o0
		);
		And270020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270000_o0,
			i1 => Or269980_o0,
			o0 => And270020_o0
		);
		Or270040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270020_o0,
			i1 => And269920_o0,
			o0 => Or270040_o0
		);
		And270060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270040_o0,
			i1 => Not1500_o0,
			o0 => And270060_o0
		);
		And270080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => And217500_o0,
			o0 => And270080_o0
		);
		And270100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270080_o0,
			i1 => Nor232220_o0,
			o0 => And270100_o0
		);
		And270120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270100_o0,
			i1 => Or219460_o0,
			o0 => And270120_o0
		);
		Or270140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270120_o0,
			i1 => And270060_o0,
			o0 => Or270140_o0
		);
		And270160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270140_o0,
			i1 => Not1080_o0,
			o0 => And270160_o0
		);
		And270180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259520_o0,
			i1 => i40,
			o0 => And270180_o0
		);
		And270200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270180_o0,
			i1 => Or267740_o0,
			o0 => And270200_o0
		);
		Or270220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270200_o0,
			i1 => And270160_o0,
			o0 => Or270220_o0
		);
		And270240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270220_o0,
			i1 => Not80_o0,
			o0 => And270240_o0
		);
		And270260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21220_o0,
			i1 => And21060_o0,
			o0 => And270260_o0
		);
		Or270280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270260_o0,
			i1 => And250120_o0,
			o0 => Or270280_o0
		);
		And270300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270280_o0,
			i1 => Not620_o0,
			o0 => And270300_o0
		);
		Or270320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270300_o0,
			i1 => And269860_o0,
			o0 => Or270320_o0
		);
		And270340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And257320_o0,
			i1 => And222800_o0,
			o0 => And270340_o0
		);
		And270360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270340_o0,
			i1 => Or270320_o0,
			o0 => And270360_o0
		);
		Or270380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270360_o0,
			i1 => And270240_o0,
			o0 => Or270380_o0
		);
		And270400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270380_o0,
			i1 => Not100_o0,
			o0 => And270400_o0
		);
		And270420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i5,
			i1 => i1,
			o0 => And270420_o0
		);
		And270440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270420_o0,
			i1 => And224500_o0,
			o0 => And270440_o0
		);
		And270460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270440_o0,
			i1 => And230760_o0,
			o0 => And270460_o0
		);
		Or270480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270460_o0,
			i1 => And270400_o0,
			o0 => Or270480_o0
		);
		And270500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270480_o0,
			i1 => Not60_o0,
			o0 => And270500_o0
		);
		And270520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And229920_o0,
			i1 => And23180_o0,
			o0 => And270520_o0
		);
		And270540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23020_o0,
			i1 => And2640_o0,
			o0 => And270540_o0
		);
		And270560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270540_o0,
			i1 => And270520_o0,
			o0 => And270560_o0
		);
		And270580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270560_o0,
			i1 => And2260_o0,
			o0 => And270580_o0
		);
		Or270600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270580_o0,
			i1 => And270500_o0,
			o0 => Or270600_o0
		);
		And270620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And220360_o0,
			i1 => And215000_o0,
			o0 => And270620_o0
		);
		And270640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270620_o0,
			i1 => Or270600_o0,
			o0 => And270640_o0
		);
		And270660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor2220_o0,
			i1 => And21300_o0,
			o0 => And270660_o0
		);
		Or270680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270660_o0,
			i1 => And28360_o0,
			o0 => Or270680_o0
		);
		And270700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270680_o0,
			i1 => i4,
			o0 => And270700_o0
		);
		And270720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28320_o0,
			i1 => Not160_o0,
			o0 => And270720_o0
		);
		Or270740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270720_o0,
			i1 => And270700_o0,
			o0 => Or270740_o0
		);
		And270760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270740_o0,
			i1 => i19,
			o0 => And270760_o0
		);
		And270780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And2640_o0,
			i1 => Not160_o0,
			o0 => And270780_o0
		);
		And270800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270780_o0,
			i1 => And269720_o0,
			o0 => And270800_o0
		);
		Or270820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270800_o0,
			i1 => And270760_o0,
			o0 => Or270820_o0
		);
		And270840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270820_o0,
			i1 => Not180_o0,
			o0 => And270840_o0
		);
		Or270860 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21640_o0,
			i1 => i15,
			o0 => Or270860_o0
		);
		Or270880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or270860_o0,
			i1 => And233100_o0,
			o0 => Or270880_o0
		);
		And270900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22100_o0,
			i1 => i40,
			o0 => And270900_o0
		);
		And270920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270900_o0,
			i1 => Or270880_o0,
			o0 => And270920_o0
		);
		Or270940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And270920_o0,
			i1 => And270840_o0,
			o0 => Or270940_o0
		);
		And270960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or270940_o0,
			i1 => i13,
			o0 => And270960_o0
		);
		And270980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor215260_o0,
			i1 => Nor21220_o0,
			o0 => And270980_o0
		);
		And271000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And270980_o0,
			i1 => And270900_o0,
			o0 => And271000_o0
		);
		And271020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271000_o0,
			i1 => Xor216780_o0,
			o0 => And271020_o0
		);
		Or271040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271020_o0,
			i1 => And270960_o0,
			o0 => Or271040_o0
		);
		And271060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271040_o0,
			i1 => Not80_o0,
			o0 => And271060_o0
		);
		And271080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22900_o0,
			i1 => And22100_o0,
			o0 => And271080_o0
		);
		And271100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271080_o0,
			i1 => And219780_o0,
			o0 => And271100_o0
		);
		And271120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271100_o0,
			i1 => And222140_o0,
			o0 => And271120_o0
		);
		Or271140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271120_o0,
			i1 => And271060_o0,
			o0 => Or271140_o0
		);
		And271160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271140_o0,
			i1 => Not540_o0,
			o0 => And271160_o0
		);
		And271180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And22400_o0,
			i1 => And21240_o0,
			o0 => And271180_o0
		);
		And271200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224500_o0,
			i1 => And215860_o0,
			o0 => And271200_o0
		);
		And271220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271200_o0,
			i1 => And271180_o0,
			o0 => And271220_o0
		);
		Or271240 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271220_o0,
			i1 => And271160_o0,
			o0 => Or271240_o0
		);
		And271260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And253960_o0,
			i1 => And23340_o0,
			o0 => And271260_o0
		);
		And271280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271260_o0,
			i1 => Or271240_o0,
			o0 => And271280_o0
		);
		Or271300 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And232660_o0,
			i1 => Not80_o0,
			o0 => Or271300_o0
		);
		And271320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271300_o0,
			i1 => i16,
			o0 => And271320_o0
		);
		Or271340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271320_o0,
			i1 => Nor252020_o0,
			o0 => Or271340_o0
		);
		And271360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And246320_o0,
			i1 => Nor23600_o0,
			o0 => And271360_o0
		);
		And271380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271360_o0,
			i1 => And253940_o0,
			o0 => And271380_o0
		);
		And271400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28140_o0,
			i1 => And23340_o0,
			o0 => And271400_o0
		);
		And271420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271400_o0,
			i1 => And271380_o0,
			o0 => And271420_o0
		);
		And271440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271420_o0,
			i1 => Or271340_o0,
			o0 => And271440_o0
		);
		And271460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And24460_o0,
			i1 => i19,
			o0 => And271460_o0
		);
		And271480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271460_o0,
			i1 => Or270680_o0,
			o0 => And271480_o0
		);
		Or271500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And28360_o0,
			i1 => i15,
			o0 => Or271500_o0
		);
		And271520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271500_o0,
			i1 => And270900_o0,
			o0 => And271520_o0
		);
		Or271540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271520_o0,
			i1 => And271480_o0,
			o0 => Or271540_o0
		);
		And271560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271540_o0,
			i1 => Not540_o0,
			o0 => And271560_o0
		);
		And271580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233000_o0,
			i1 => And215860_o0,
			o0 => And271580_o0
		);
		And271600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271580_o0,
			i1 => And270260_o0,
			o0 => And271600_o0
		);
		Or271620 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271600_o0,
			i1 => And271560_o0,
			o0 => Or271620_o0
		);
		And271640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => Nor23280_o0,
			o0 => And271640_o0
		);
		And271660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271640_o0,
			i1 => And28160_o0,
			o0 => And271660_o0
		);
		And271680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271660_o0,
			i1 => And23340_o0,
			o0 => And271680_o0
		);
		And271700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271680_o0,
			i1 => Or271620_o0,
			o0 => And271700_o0
		);
		And271720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => Not160_o0,
			o0 => And271720_o0
		);
		And271740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271720_o0,
			i1 => And215440_o0,
			o0 => And271740_o0
		);
		Or271760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271740_o0,
			i1 => And270700_o0,
			o0 => Or271760_o0
		);
		And271780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271760_o0,
			i1 => i19,
			o0 => And271780_o0
		);
		And271800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21300_o0,
			i1 => Not160_o0,
			o0 => And271800_o0
		);
		And271820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And271800_o0,
			i1 => And269720_o0,
			o0 => And271820_o0
		);
		Or271840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271820_o0,
			i1 => And271780_o0,
			o0 => Or271840_o0
		);
		And271860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271840_o0,
			i1 => Not180_o0,
			o0 => And271860_o0
		);
		Or271880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And233100_o0,
			i1 => i15,
			o0 => Or271880_o0
		);
		And271900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271880_o0,
			i1 => And270900_o0,
			o0 => And271900_o0
		);
		Or271920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271900_o0,
			i1 => And271860_o0,
			o0 => Or271920_o0
		);
		And271940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271920_o0,
			i1 => Not80_o0,
			o0 => And271940_o0
		);
		And271960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255140_o0,
			i1 => And22100_o0,
			o0 => And271960_o0
		);
		Or271980 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And271960_o0,
			i1 => And271940_o0,
			o0 => Or271980_o0
		);
		And272000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or271980_o0,
			i1 => Not540_o0,
			o0 => And272000_o0
		);
		And272020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215860_o0,
			i1 => Nor24000_o0,
			o0 => And272020_o0
		);
		And272040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272020_o0,
			i1 => And271180_o0,
			o0 => And272040_o0
		);
		Or272060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272040_o0,
			i1 => And272000_o0,
			o0 => Or272060_o0
		);
		And272080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272060_o0,
			i1 => i13,
			o0 => And272080_o0
		);
		And272100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And260480_o0,
			i1 => And215860_o0,
			o0 => And272100_o0
		);
		And272120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272100_o0,
			i1 => And23060_o0,
			o0 => And272120_o0
		);
		Or272140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272120_o0,
			i1 => And272080_o0,
			o0 => Or272140_o0
		);
		And272160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272140_o0,
			i1 => And271260_o0,
			o0 => And272160_o0
		);
		And272180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And225320_o0,
			i1 => And28040_o0,
			o0 => And272180_o0
		);
		And272200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272180_o0,
			i1 => Nor232220_o0,
			o0 => And272200_o0
		);
		And272220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272200_o0,
			i1 => Not7440_o0,
			o0 => And272220_o0
		);
		And272240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => i5,
			o0 => And272240_o0
		);
		And272260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272240_o0,
			i1 => And226440_o0,
			o0 => And272260_o0
		);
		Or272280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272260_o0,
			i1 => And272220_o0,
			o0 => Or272280_o0
		);
		Nor272300 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i18,
			o0 => Nor272300_o0
		);
		And272320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor272300_o0,
			i1 => Nor212640_o0,
			o0 => And272320_o0
		);
		And272340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor220340_o0,
			i1 => Nor214960_o0,
			o0 => And272340_o0
		);
		And272360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272340_o0,
			i1 => And28160_o0,
			o0 => And272360_o0
		);
		And272380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272360_o0,
			i1 => And272320_o0,
			o0 => And272380_o0
		);
		And272400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272380_o0,
			i1 => Or272280_o0,
			o0 => And272400_o0
		);
		Or272420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And21060_o0,
			i1 => Not80_o0,
			o0 => Or272420_o0
		);
		And272440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272420_o0,
			i1 => And271420_o0,
			o0 => And272440_o0
		);
		And272460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor226020_o0,
			i1 => Nor212700_o0,
			o0 => And272460_o0
		);
		And272480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272460_o0,
			i1 => And227400_o0,
			o0 => And272480_o0
		);
		Nor272500 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i36,
			i1 => i19,
			o0 => Nor272500_o0
		);
		And272520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor272500_o0,
			i1 => And210100_o0,
			o0 => And272520_o0
		);
		And272540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272520_o0,
			i1 => And228980_o0,
			o0 => And272540_o0
		);
		And272560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272540_o0,
			i1 => And272480_o0,
			o0 => And272560_o0
		);
		And272580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272560_o0,
			i1 => And240040_o0,
			o0 => And272580_o0
		);
		And272600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And249020_o0,
			i1 => And213280_o0,
			o0 => And272600_o0
		);
		And272620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228580_o0,
			i1 => Not80_o0,
			o0 => And272620_o0
		);
		And272640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272620_o0,
			i1 => And259520_o0,
			o0 => And272640_o0
		);
		And272660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219520_o0,
			i1 => Nor264380_o0,
			o0 => And272660_o0
		);
		Or272680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272660_o0,
			i1 => And272640_o0,
			o0 => Or272680_o0
		);
		And272700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272680_o0,
			i1 => Not180_o0,
			o0 => And272700_o0
		);
		And272720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => And22300_o0,
			o0 => And272720_o0
		);
		Or272740 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272720_o0,
			i1 => And219920_o0,
			o0 => Or272740_o0
		);
		And272760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272740_o0,
			i1 => And211020_o0,
			o0 => And272760_o0
		);
		Or272780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272760_o0,
			i1 => And272700_o0,
			o0 => Or272780_o0
		);
		And272800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272780_o0,
			i1 => i16,
			o0 => And272800_o0
		);
		And272820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i5,
			o0 => And272820_o0
		);
		And272840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272820_o0,
			i1 => And22300_o0,
			o0 => And272840_o0
		);
		Nor272860 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i14,
			i1 => i5,
			o0 => Nor272860_o0
		);
		And272880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And28060_o0,
			i1 => i5,
			o0 => And272880_o0
		);
		Or272900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272880_o0,
			i1 => Nor272860_o0,
			o0 => Or272900_o0
		);
		Or272920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or272900_o0,
			i1 => And272840_o0,
			o0 => Or272920_o0
		);
		And272940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or272920_o0,
			i1 => Nor224000_o0,
			o0 => And272940_o0
		);
		And272960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And228580_o0,
			i1 => i14,
			o0 => And272960_o0
		);
		And272980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And272960_o0,
			i1 => And250340_o0,
			o0 => And272980_o0
		);
		And273000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor232220_o0,
			i1 => And219900_o0,
			o0 => And273000_o0
		);
		And273020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And213180_o0,
			i1 => And211020_o0,
			o0 => And273020_o0
		);
		Or273040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273020_o0,
			i1 => And273000_o0,
			o0 => Or273040_o0
		);
		And273060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And212880_o0,
			i1 => And22480_o0,
			o0 => And273060_o0
		);
		And273080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273060_o0,
			i1 => Or273040_o0,
			o0 => And273080_o0
		);
		Or273100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273080_o0,
			i1 => And272980_o0,
			o0 => Or273100_o0
		);
		Or273120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or273100_o0,
			i1 => And272940_o0,
			o0 => Or273120_o0
		);
		Or273140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or273120_o0,
			i1 => And272800_o0,
			o0 => Or273140_o0
		);
		And273160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or273140_o0,
			i1 => And26520_o0,
			o0 => And273160_o0
		);
		And273180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And227520_o0,
			i1 => And23020_o0,
			o0 => And273180_o0
		);
		And273200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273180_o0,
			i1 => And224180_o0,
			o0 => And273200_o0
		);
		Or273220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273200_o0,
			i1 => And273160_o0,
			o0 => Or273220_o0
		);
		And273240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And259520_o0,
			i1 => And213180_o0,
			o0 => And273240_o0
		);
		And273260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273240_o0,
			i1 => And21960_o0,
			o0 => And273260_o0
		);
		Or273280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273260_o0,
			i1 => And220160_o0,
			o0 => Or273280_o0
		);
		And273300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or273280_o0,
			i1 => i12,
			o0 => And273300_o0
		);
		And273320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And223260_o0,
			i1 => Nor21840_o0,
			o0 => And273320_o0
		);
		And273340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273320_o0,
			i1 => Nor232220_o0,
			o0 => And273340_o0
		);
		And273360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273340_o0,
			i1 => And21240_o0,
			o0 => And273360_o0
		);
		Or273380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273360_o0,
			i1 => And273300_o0,
			o0 => Or273380_o0
		);
		And273400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or273380_o0,
			i1 => And26520_o0,
			o0 => And273400_o0
		);
		Or273420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273400_o0,
			i1 => Or273220_o0,
			o0 => Or273420_o0
		);
		And273440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or273420_o0,
			i1 => Not12100_o0,
			o0 => And273440_o0
		);
		And273460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor240760_o0,
			i1 => i8,
			o0 => And273460_o0
		);
		Or273480 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273460_o0,
			i1 => And273440_o0,
			o0 => Or273480_o0
		);
		And273500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or273480_o0,
			i1 => Not24960_o0,
			o0 => And273500_o0
		);
		And273520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i11,
			i1 => i8,
			o0 => And273520_o0
		);
		And273540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273520_o0,
			i1 => Nor240760_o0,
			o0 => And273540_o0
		);
		Or273560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273540_o0,
			i1 => And273500_o0,
			o0 => Or273560_o0
		);
		And273580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or273560_o0,
			i1 => Not12120_o0,
			o0 => And273580_o0
		);
		And273600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i10,
			i1 => i8,
			o0 => And273600_o0
		);
		And273620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273600_o0,
			i1 => Nor240760_o0,
			o0 => And273620_o0
		);
		Or273640 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273620_o0,
			i1 => And273580_o0,
			o0 => Or273640_o0
		);
		And273660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263280_o0,
			i1 => Nor226140_o0,
			o0 => And273660_o0
		);
		And273680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273660_o0,
			i1 => Or273640_o0,
			o0 => And273680_o0
		);
		Or273700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And228840_o0,
			i1 => And226520_o0,
			o0 => Or273700_o0
		);
		And273720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23080_o0,
			i1 => Not1080_o0,
			o0 => And273720_o0
		);
		And273740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273720_o0,
			i1 => Or273700_o0,
			o0 => And273740_o0
		);
		Nor273760 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => Not1080_o0,
			o0 => Nor273760_o0
		);
		And273780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor273760_o0,
			i1 => And22800_o0,
			o0 => And273780_o0
		);
		And273800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273780_o0,
			i1 => And23020_o0,
			o0 => And273800_o0
		);
		Or273820 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273800_o0,
			i1 => And273740_o0,
			o0 => Or273820_o0
		);
		And273840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216820_o0,
			i1 => And25600_o0,
			o0 => And273840_o0
		);
		And273860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214960_o0,
			i1 => Nor212640_o0,
			o0 => And273860_o0
		);
		And273880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273860_o0,
			i1 => And273840_o0,
			o0 => And273880_o0
		);
		And273900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273880_o0,
			i1 => Or273820_o0,
			o0 => And273900_o0
		);
		Or273920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And273900_o0,
			i1 => i8,
			o0 => Or273920_o0
		);
		And273940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263280_o0,
			i1 => And23620_o0,
			o0 => And273940_o0
		);
		And273960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273940_o0,
			i1 => Or273920_o0,
			o0 => And273960_o0
		);
		Nor273980 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i38,
			i1 => i37,
			o0 => Nor273980_o0
		);
		Nor274000 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i36,
			o0 => Nor274000_o0
		);
		And274020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor274000_o0,
			i1 => Nor273980_o0,
			o0 => And274020_o0
		);
		And274040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => And212880_o0,
			o0 => And274040_o0
		);
		And274060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23520_o0,
			i1 => And21300_o0,
			o0 => And274060_o0
		);
		And274080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274060_o0,
			i1 => And274040_o0,
			o0 => And274080_o0
		);
		And274100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274080_o0,
			i1 => And274020_o0,
			o0 => And274100_o0
		);
		And274120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255560_o0,
			i1 => Nor232220_o0,
			o0 => And274120_o0
		);
		And274140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274120_o0,
			i1 => And240040_o0,
			o0 => And274140_o0
		);
		And274160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274140_o0,
			i1 => And274100_o0,
			o0 => And274160_o0
		);
		Or274180 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And244220_o0,
			i1 => i14,
			o0 => Or274180_o0
		);
		And274200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274180_o0,
			i1 => And211940_o0,
			o0 => And274200_o0
		);
		And274220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not1280_o0,
			i1 => i14,
			o0 => And274220_o0
		);
		And274240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274220_o0,
			i1 => And214100_o0,
			o0 => And274240_o0
		);
		And274260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219620_o0,
			i1 => Nor214120_o0,
			o0 => And274260_o0
		);
		Or274280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274260_o0,
			i1 => And274240_o0,
			o0 => Or274280_o0
		);
		And274300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274280_o0,
			i1 => i13,
			o0 => And274300_o0
		);
		And274320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => i17,
			o0 => And274320_o0
		);
		And274340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274320_o0,
			i1 => Not7440_o0,
			o0 => And274340_o0
		);
		Or274360 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274340_o0,
			i1 => And274300_o0,
			o0 => Or274360_o0
		);
		And274380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274360_o0,
			i1 => Not1080_o0,
			o0 => And274380_o0
		);
		And274400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor252020_o0,
			i1 => And2260_o0,
			o0 => And274400_o0
		);
		Or274420 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274400_o0,
			i1 => i14,
			o0 => Or274420_o0
		);
		And274440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274420_o0,
			i1 => Not2080_o0,
			o0 => And274440_o0
		);
		Or274460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274440_o0,
			i1 => And274380_o0,
			o0 => Or274460_o0
		);
		And274480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274460_o0,
			i1 => Not620_o0,
			o0 => And274480_o0
		);
		And274500 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => And23780_o0,
			o0 => And274500_o0
		);
		And274520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And263580_o0,
			i1 => And234780_o0,
			o0 => And274520_o0
		);
		Or274540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274520_o0,
			i1 => And274500_o0,
			o0 => Or274540_o0
		);
		Or274560 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or274540_o0,
			i1 => And274480_o0,
			o0 => Or274560_o0
		);
		Or274580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or274560_o0,
			i1 => And274200_o0,
			o0 => Or274580_o0
		);
		And274600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274580_o0,
			i1 => i12,
			o0 => And274600_o0
		);
		And274620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And21940_o0,
			i1 => And21100_o0,
			o0 => And274620_o0
		);
		And274640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219900_o0,
			i1 => And23020_o0,
			o0 => And274640_o0
		);
		And274660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274640_o0,
			i1 => And274620_o0,
			o0 => And274660_o0
		);
		Or274680 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274660_o0,
			i1 => And274600_o0,
			o0 => Or274680_o0
		);
		And274700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274680_o0,
			i1 => And26520_o0,
			o0 => And274700_o0
		);
		Or274720 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274700_o0,
			i1 => And257980_o0,
			o0 => Or274720_o0
		);
		And274740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274720_o0,
			i1 => Not60_o0,
			o0 => And274740_o0
		);
		Or274760 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274740_o0,
			i1 => And264980_o0,
			o0 => Or274760_o0
		);
		And274780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274760_o0,
			i1 => And265040_o0,
			o0 => And274780_o0
		);
		And274800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or261840_o0,
			i1 => Or210400_o0,
			o0 => And274800_o0
		);
		And274820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => i26,
			o0 => And274820_o0
		);
		And274840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274820_o0,
			i1 => And254820_o0,
			o0 => And274840_o0
		);
		And274860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And234540_o0,
			i1 => Nor234140_o0,
			o0 => And274860_o0
		);
		And274880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274860_o0,
			i1 => And274840_o0,
			o0 => And274880_o0
		);
		Or274900 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And274880_o0,
			i1 => And274800_o0,
			o0 => Or274900_o0
		);
		And274920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or274900_o0,
			i1 => Nor226140_o0,
			o0 => And274920_o0
		);
		Xor274940 : entity gtech_lib.xor2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => i2,
			o0 => Xor274940_o0
		);
		And274960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Xor274940_o0,
			i1 => And210540_o0,
			o0 => And274960_o0
		);
		And274980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i4,
			i1 => Not120_o0,
			o0 => And274980_o0
		);
		And275000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And274980_o0,
			i1 => And210600_o0,
			o0 => And275000_o0
		);
		Or275020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275000_o0,
			i1 => And274960_o0,
			o0 => Or275020_o0
		);
		Or275040 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => Or275020_o0,
			i1 => And274920_o0,
			o0 => Or275040_o0
		);
		And275060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275040_o0,
			i1 => i27,
			o0 => And275060_o0
		);
		And275080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or210620_o0,
			i1 => Or210400_o0,
			o0 => And275080_o0
		);
		Or275100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => i24,
			i1 => i23,
			o0 => Or275100_o0
		);
		And275120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275100_o0,
			i1 => i22,
			o0 => And275120_o0
		);
		Or275140 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275120_o0,
			i1 => And210740_o0,
			o0 => Or275140_o0
		);
		And275160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And261940_o0,
			i1 => Nor234140_o0,
			o0 => And275160_o0
		);
		And275180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275160_o0,
			i1 => Or275140_o0,
			o0 => And275180_o0
		);
		Or275200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275180_o0,
			i1 => And275080_o0,
			o0 => Or275200_o0
		);
		And275220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275200_o0,
			i1 => Not9580_o0,
			o0 => And275220_o0
		);
		And275240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i20,
			i1 => Not540_o0,
			o0 => And275240_o0
		);
		And275260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275240_o0,
			i1 => And261940_o0,
			o0 => And275260_o0
		);
		Or275280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275260_o0,
			i1 => And275220_o0,
			o0 => Or275280_o0
		);
		And275300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275280_o0,
			i1 => Nor226140_o0,
			o0 => And275300_o0
		);
		Or275320 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275300_o0,
			i1 => And275060_o0,
			o0 => Or275320_o0
		);
		And275340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275320_o0,
			i1 => Not1500_o0,
			o0 => And275340_o0
		);
		And275360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor226140_o0,
			i1 => Not540_o0,
			o0 => And275360_o0
		);
		And275380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275360_o0,
			i1 => And224580_o0,
			o0 => And275380_o0
		);
		Or275400 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275380_o0,
			i1 => And275340_o0,
			o0 => Or275400_o0
		);
		And275420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275400_o0,
			i1 => And26580_o0,
			o0 => And275420_o0
		);
		And275440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not120_o0,
			o0 => And275440_o0
		);
		And275460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And224580_o0,
			i1 => And24620_o0,
			o0 => And275460_o0
		);
		And275480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275460_o0,
			i1 => And275440_o0,
			o0 => And275480_o0
		);
		Or275500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275480_o0,
			i1 => And275420_o0,
			o0 => Or275500_o0
		);
		And275520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275500_o0,
			i1 => Not140_o0,
			o0 => And275520_o0
		);
		And275540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And215860_o0,
			i1 => And26040_o0,
			o0 => And275540_o0
		);
		And275560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275540_o0,
			i1 => And254620_o0,
			o0 => And275560_o0
		);
		And275580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275560_o0,
			i1 => And218280_o0,
			o0 => And275580_o0
		);
		Or275600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275580_o0,
			i1 => And275520_o0,
			o0 => Or275600_o0
		);
		And275620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not3300_o0,
			i1 => i17,
			o0 => And275620_o0
		);
		And275640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275620_o0,
			i1 => Nor24920_o0,
			o0 => And275640_o0
		);
		And275660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor23320_o0,
			i1 => And23080_o0,
			o0 => And275660_o0
		);
		And275680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275660_o0,
			i1 => And256660_o0,
			o0 => And275680_o0
		);
		And275700 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275680_o0,
			i1 => And275640_o0,
			o0 => And275700_o0
		);
		And275720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275700_o0,
			i1 => Or275600_o0,
			o0 => And275720_o0
		);
		Nor275740 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => Xor218020_o0,
			i1 => Not540_o0,
			o0 => Nor275740_o0
		);
		And275760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And29720_o0,
			i1 => Not540_o0,
			o0 => And275760_o0
		);
		Or275780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275760_o0,
			i1 => Nor275740_o0,
			o0 => Or275780_o0
		);
		And275800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275780_o0,
			i1 => And26040_o0,
			o0 => And275800_o0
		);
		And275820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And255620_o0,
			i1 => And221240_o0,
			o0 => And275820_o0
		);
		Or275840 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275820_o0,
			i1 => And275800_o0,
			o0 => Or275840_o0
		);
		And275860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275840_o0,
			i1 => Not160_o0,
			o0 => And275860_o0
		);
		And275880 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221240_o0,
			i1 => i5,
			o0 => And275880_o0
		);
		And275900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275880_o0,
			i1 => And238720_o0,
			o0 => And275900_o0
		);
		Or275920 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And275900_o0,
			i1 => And275860_o0,
			o0 => Or275920_o0
		);
		And275940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or275920_o0,
			i1 => Nand210560_o0,
			o0 => And275940_o0
		);
		And275960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or217820_o0,
			i1 => i4,
			o0 => And275960_o0
		);
		And275980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i22,
			i1 => Not160_o0,
			o0 => And275980_o0
		);
		And276000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And275980_o0,
			i1 => And263020_o0,
			o0 => And276000_o0
		);
		Or276020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276000_o0,
			i1 => And275960_o0,
			o0 => Or276020_o0
		);
		And276040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276020_o0,
			i1 => i27,
			o0 => And276040_o0
		);
		And276060 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Not9580_o0,
			i1 => i23,
			o0 => And276060_o0
		);
		And276080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276060_o0,
			i1 => And275980_o0,
			o0 => And276080_o0
		);
		Or276100 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276080_o0,
			i1 => And276040_o0,
			o0 => Or276100_o0
		);
		And276120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276100_o0,
			i1 => Not540_o0,
			o0 => And276120_o0
		);
		And276140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And221280_o0,
			i1 => And215860_o0,
			o0 => And276140_o0
		);
		Or276160 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276140_o0,
			i1 => And276120_o0,
			o0 => Or276160_o0
		);
		And276180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276160_o0,
			i1 => And26040_o0,
			o0 => And276180_o0
		);
		Or276200 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276180_o0,
			i1 => And275940_o0,
			o0 => Or276200_o0
		);
		And276220 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276200_o0,
			i1 => And238360_o0,
			o0 => And276220_o0
		);
		And276240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor235820_o0,
			i1 => Nor22600_o0,
			o0 => And276240_o0
		);
		And276260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276240_o0,
			i1 => And24940_o0,
			o0 => And276260_o0
		);
		Or276280 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276260_o0,
			i1 => And276220_o0,
			o0 => Or276280_o0
		);
		And276300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And23700_o0,
			i1 => Nor23600_o0,
			o0 => And276300_o0
		);
		And276320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor272500_o0,
			i1 => And21940_o0,
			o0 => And276320_o0
		);
		And276340 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => And23080_o0,
			o0 => And276340_o0
		);
		And276360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276340_o0,
			i1 => And276320_o0,
			o0 => And276360_o0
		);
		And276380 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276360_o0,
			i1 => And276300_o0,
			o0 => And276380_o0
		);
		And276400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276380_o0,
			i1 => Or276280_o0,
			o0 => And276400_o0
		);
		And276420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And219600_o0,
			i1 => Not1040_o0,
			o0 => And276420_o0
		);
		Or276440 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276420_o0,
			i1 => And29280_o0,
			o0 => Or276440_o0
		);
		And276460 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276440_o0,
			i1 => i15,
			o0 => And276460_o0
		);
		And276480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And231420_o0,
			i1 => Nor29260_o0,
			o0 => And276480_o0
		);
		Or276500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276480_o0,
			i1 => And276460_o0,
			o0 => Or276500_o0
		);
		And276520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276500_o0,
			i1 => And2560_o0,
			o0 => And276520_o0
		);
		And276540 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor24920_o0,
			i1 => i17,
			o0 => And276540_o0
		);
		And276560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276540_o0,
			i1 => And219500_o0,
			o0 => And276560_o0
		);
		And276580 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276560_o0,
			i1 => And215220_o0,
			o0 => And276580_o0
		);
		Or276600 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276580_o0,
			i1 => And276520_o0,
			o0 => Or276600_o0
		);
		And276620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276600_o0,
			i1 => Not160_o0,
			o0 => And276620_o0
		);
		And276640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor211040_o0,
			i1 => i17,
			o0 => And276640_o0
		);
		And276660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276640_o0,
			i1 => And230240_o0,
			o0 => And276660_o0
		);
		And276680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276660_o0,
			i1 => And211200_o0,
			o0 => And276680_o0
		);
		Or276700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276680_o0,
			i1 => And276620_o0,
			o0 => Or276700_o0
		);
		And276720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276700_o0,
			i1 => i18,
			o0 => And276720_o0
		);
		And276740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => Nor21260_o0,
			o0 => And276740_o0
		);
		And276760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276740_o0,
			i1 => And228580_o0,
			o0 => And276760_o0
		);
		And276780 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276760_o0,
			i1 => And224600_o0,
			o0 => And276780_o0
		);
		Or276800 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276780_o0,
			i1 => And276720_o0,
			o0 => Or276800_o0
		);
		And276820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276800_o0,
			i1 => Not1280_o0,
			o0 => And276820_o0
		);
		And276840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216160_o0,
			i1 => i16,
			o0 => And276840_o0
		);
		And276860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276840_o0,
			i1 => Nor24920_o0,
			o0 => And276860_o0
		);
		Or276880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276860_o0,
			i1 => And28060_o0,
			o0 => Or276880_o0
		);
		And276900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not2080_o0,
			o0 => And276900_o0
		);
		And276920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276900_o0,
			i1 => Nor21260_o0,
			o0 => And276920_o0
		);
		And276940 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And276920_o0,
			i1 => Or276880_o0,
			o0 => And276940_o0
		);
		Or276960 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And276940_o0,
			i1 => And276820_o0,
			o0 => Or276960_o0
		);
		And276980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or276960_o0,
			i1 => Not60_o0,
			o0 => And276980_o0
		);
		And277000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => Not540_o0,
			o0 => And277000_o0
		);
		And277020 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277000_o0,
			i1 => And214620_o0,
			o0 => And277020_o0
		);
		And277040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277020_o0,
			i1 => And23060_o0,
			o0 => And277040_o0
		);
		Or277060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277040_o0,
			i1 => And276980_o0,
			o0 => Or277060_o0
		);
		And277080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214980_o0,
			i1 => i12,
			o0 => And277080_o0
		);
		And277100 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor214960_o0,
			i1 => Nor214740_o0,
			o0 => And277100_o0
		);
		And277120 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277100_o0,
			i1 => Nor22060_o0,
			o0 => And277120_o0
		);
		And277140 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277120_o0,
			i1 => And277080_o0,
			o0 => And277140_o0
		);
		And277160 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277140_o0,
			i1 => Or277060_o0,
			o0 => And277160_o0
		);
		And277180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i16,
			i1 => i14,
			o0 => And277180_o0
		);
		And277200 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277180_o0,
			i1 => Nor214120_o0,
			o0 => And277200_o0
		);
		Or277220 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277200_o0,
			i1 => Nor252020_o0,
			o0 => Or277220_o0
		);
		And277240 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277220_o0,
			i1 => And271420_o0,
			o0 => And277240_o0
		);
		And277260 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And269860_o0,
			i1 => And219600_o0,
			o0 => And277260_o0
		);
		And277280 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor29260_o0,
			i1 => Nor21840_o0,
			o0 => And277280_o0
		);
		And277300 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And216820_o0,
			i1 => And210100_o0,
			o0 => And277300_o0
		);
		And277320 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277300_o0,
			i1 => And277280_o0,
			o0 => And277320_o0
		);
		Or277340 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277320_o0,
			i1 => And277260_o0,
			o0 => Or277340_o0
		);
		And277360 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277340_o0,
			i1 => Not540_o0,
			o0 => And277360_o0
		);
		Or277380 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277360_o0,
			i1 => And220020_o0,
			o0 => Or277380_o0
		);
		And277400 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277380_o0,
			i1 => i19,
			o0 => And277400_o0
		);
		And277420 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21840_o0,
			i1 => i14,
			o0 => And277420_o0
		);
		And277440 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277420_o0,
			i1 => And21820_o0,
			o0 => And277440_o0
		);
		Or277460 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277440_o0,
			i1 => And226800_o0,
			o0 => Or277460_o0
		);
		And277480 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277460_o0,
			i1 => And259520_o0,
			o0 => And277480_o0
		);
		Or277500 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277480_o0,
			i1 => And277400_o0,
			o0 => Or277500_o0
		);
		And277520 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277500_o0,
			i1 => i12,
			o0 => And277520_o0
		);
		Or277540 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277520_o0,
			i1 => And273360_o0,
			o0 => Or277540_o0
		);
		And277560 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277540_o0,
			i1 => And26520_o0,
			o0 => And277560_o0
		);
		Or277580 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277560_o0,
			i1 => Or273220_o0,
			o0 => Or277580_o0
		);
		And277600 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And256660_o0,
			i1 => Nor226140_o0,
			o0 => And277600_o0
		);
		And277620 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277600_o0,
			i1 => And23340_o0,
			o0 => And277620_o0
		);
		And277640 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277620_o0,
			i1 => Or277580_o0,
			o0 => And277640_o0
		);
		And277660 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And273720_o0,
			i1 => Or220780_o0,
			o0 => And277660_o0
		);
		And277680 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And233660_o0,
			i1 => And212900_o0,
			o0 => And277680_o0
		);
		Or277700 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277680_o0,
			i1 => And277660_o0,
			o0 => Or277700_o0
		);
		And277720 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277700_o0,
			i1 => Not1500_o0,
			o0 => And277720_o0
		);
		And277740 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor22900_o0,
			i1 => And2240_o0,
			o0 => And277740_o0
		);
		And277760 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277740_o0,
			i1 => And233660_o0,
			o0 => And277760_o0
		);
		Or277780 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277760_o0,
			i1 => And277720_o0,
			o0 => Or277780_o0
		);
		And277800 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or277780_o0,
			i1 => Not20760_o0,
			o0 => And277800_o0
		);
		And277820 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i39,
			i1 => i19,
			o0 => And277820_o0
		);
		And277840 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277820_o0,
			i1 => And210100_o0,
			o0 => And277840_o0
		);
		And277860 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277840_o0,
			i1 => And230540_o0,
			o0 => And277860_o0
		);
		Or277880 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277860_o0,
			i1 => And277800_o0,
			o0 => Or277880_o0
		);
		And277900 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => i40,
			i1 => Not80_o0,
			o0 => And277900_o0
		);
		And277920 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277900_o0,
			i1 => Or277880_o0,
			o0 => And277920_o0
		);
		Or277940 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And277920_o0,
			i1 => Not24560_o0,
			o0 => Or277940_o0
		);
		And277960 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor21260_o0,
			i1 => Not3300_o0,
			o0 => And277960_o0
		);
		And277980 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277960_o0,
			i1 => And28160_o0,
			o0 => And277980_o0
		);
		And278000 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => And277980_o0,
			i1 => Or277940_o0,
			o0 => And278000_o0
		);
		Or278020 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And278000_o0,
			i1 => i36,
			o0 => Or278020_o0
		);
		And278040 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or278020_o0,
			i1 => Nor212700_o0,
			o0 => And278040_o0
		);
		Or278060 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And278040_o0,
			i1 => And220740_o0,
			o0 => Or278060_o0
		);
		And278080 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Or278060_o0,
			i1 => Nor255540_o0,
			o0 => And278080_o0
		);
		Or279120 : entity gtech_lib.or2_d
		generic map(1000 fs)
		port map(
			i0 => And272580_o0,
			i1 => And279180_o0,
			o0 => Or279120_o0
		);
		Nor279140 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => And268860_o0,
			i1 => And25800_o0,
			o0 => Nor279140_o0
		);
		Nor279160 : entity gtech_lib.nor2_d
		generic map(1000 fs)
		port map(
			i0 => And245140_o0,
			i1 => Nand210020_o0,
			o0 => Nor279160_o0
		);
		And279180 : entity gtech_lib.and2_d
		generic map(1000 fs)
		port map(
			i0 => Nor279140_o0,
			i1 => Nor279160_o0,
			o0 => And279180_o0
		);
	----------------------------------
	-- Wiring primary ouputs 
	----------------------------------
	o0 <= And23380_o0;
	o1 <= '0';
	o2 <= And23760_o0;
	o3 <= And23960_o0;
	o4 <= And26960_o0;
	o5 <= And28240_o0;
	o6 <= And29400_o0;
	o7 <= And212080_o0;
	o8 <= And212820_o0;
	o9 <= And213320_o0;
	o10 <= And213640_o0;
	o11 <= And214840_o0;
	o12 <= And215040_o0;
	o13 <= And215800_o0;
	o14 <= And219160_o0;
	o15 <= Or220720_o0;
	o16 <= And225040_o0;
	o17 <= And225440_o0;
	o18 <= Or226300_o0;
	o19 <= Or227700_o0;
	o20 <= And231200_o0;
	o21 <= And231380_o0;
	o22 <= Or235100_o0;
	o23 <= And235360_o0;
	o24 <= Or240240_o0;
	o25 <= And242240_o0;
	o26 <= And244780_o0;
	o27 <= Or248960_o0;
	o28 <= And249120_o0;
	o29 <= Or251060_o0;
	o30 <= And251160_o0;
	o31 <= '0';
	o32 <= '0';
	o33 <= And251220_o0;
	o34 <= Or251840_o0;
	o35 <= And251900_o0;
	o36 <= And252180_o0;
	o37 <= Or253080_o0;
	o38 <= Or253820_o0;
	o39 <= '0';
	o40 <= And254040_o0;
	o41 <= And255600_o0;
	o42 <= And256700_o0;
	o43 <= And258180_o0;
	o44 <= And259300_o0;
	o45 <= And260600_o0;
	o46 <= And261760_o0;
	o47 <= And263440_o0;
	o48 <= And265060_o0;
	o49 <= And265680_o0;
	o50 <= And267080_o0;
	o51 <= And268660_o0;
	o52 <= And269820_o0;
	o53 <= And270640_o0;
	o54 <= And271280_o0;
	o55 <= And271440_o0;
	o56 <= And271700_o0;
	o57 <= And272160_o0;
	o58 <= And272400_o0;
	o59 <= And272440_o0;
	o60 <= Or279120_o0;
	o61 <= And272600_o0;
	o62 <= And273680_o0;
	o63 <= And273960_o0;
	o64 <= And274160_o0;
	o65 <= And274780_o0;
	o66 <= And275720_o0;
	o67 <= And276400_o0;
	o68 <= And277160_o0;
	o69 <= And277240_o0;
	o70 <= And277640_o0;
	o71 <= And220680_o0;
	o72 <= And278080_o0;
end netenos;
